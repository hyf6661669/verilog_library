接"test_0.sv"测试一下Radix-4 SRT计算整数除法时余数的求法.
在"test_2.sv"中有更精确的描述, 这部分内容不用看了. 先保留着不删了吧。

// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 001111111111001010100011 = 4190883
D[24-1:0] = 000000000010101011110001 = 10993
Q[24-1:0] = X / D = 381 = 000000000000000101111101
REM[24-1:0] = 4190883 - 381 * 10993 = 2550 = 000000000000100111110110
按照小数除法的方式, 将X和D规格化:
CLZ_X = 2
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 8
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 5
Dividend[25-1:0] 	= 0_111111111100101010001100
Divisor[25-1:0] 	= 0_101010111100010000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -16 	= 111_0000
m[0] 	= -6 	= 111_1001
m[1] 	= 4		= 000_0100
m[2] 	= 15	= 000_1111

+ D = 000_10101011110001000000000000
+2D = 001_01010111100010000000000000
- D = 111_01010100001111000000000000
-2D = 110_10101000011110000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[5] = 0_00100111110110000000000000 >= 0
q[final] = q[5]
q_pos = 1000_0000_01
q_neg = 0010_0001_00
q_calculated_pre = q_pos - q_neg = 0101111101
q_calculated = q_calculated_pre - (w[final] < 0) = 0101111101
remainder[24-1:0] = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
001001111101100000000000 >> 10 = 
000000000000100111110110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00111111111100101010001100
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[2], +Inf)" -> q[1] = +2
q_pos = 10
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_11111111110010101000110000 + 
110_10101000011110000000000000 = 
111_10101000010000101000110000 -> 
w[1] = 1_10101000010000101000110000
4 * w[1] = 110_10100001000010100011000000
(4 * w[1])_trunc_3_4 = 110_1010, "belongs to [-Inf, m[-1])" -> q[2] = -2
q_pos = 1000
q_neg = 0010

ITER[1]:
4 * w[1] + (-q[2] * D) = 
110_10100001000010100011000000 + 
001_01010111100010000000000000 = 
111_11111000100100100011000000 -> 
w[2] = 1_11111000100100100011000000
4 * w[2] = 111_11100010010010001100000000
(4 * w[2])_trunc_3_4 = 111_1110, "belongs to [m[0], m[1])" -> q[3] = 0
q_pos = 1000_00
q_neg = 0010_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_11100010010010001100000000 + 
000_00000000000000000000000000 = 
111_11100010010010001100000000 -> 
w[3] = 1_11100010010010001100000000
4 * w[3] = 111_10001001001000110000000000
(4 * w[3])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 1000_0000
q_neg = 0010_0001

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_10001001001000110000000000 + 
000_10101011110001000000000000 = 
000_00110100111001110000000000 -> 
w[4] = 0_00110100111001110000000000
4 * w[4] = 000_11010011100111000000000000
(4 * w[4])_trunc_3_4 = 000_0101, "belongs to [m[1], m[2])" -> q[5] = +1
q_pos = 1000_0000_01
q_neg = 0010_0001_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
000_11010011100111000000000000 + 
111_01010100001111000000000000 = 
000_00100111110110000000000000 -> 
w[5] = 0_00100111110110000000000000
4 * w[5] = 000_10011111011000000000000000
(4 * w[5])_trunc_3_4 = 000_1001, "belongs to [m[1], m[2])" -> q[6] = +1
q_pos = 1000_0000_0101
q_neg = 0010_0001_0000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 000000000000000001111101 = 125
D[24-1:0] = 000000000000000000000110 = 6

CLZ_X = 17
CLZ_D = 21
CLZ_DIFF = CLZ_D - CLZ_X = 4
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 3
Dividend[25-1:0] 	= 0_111110100000000000000000
Divisor[25-1:0] 	= 0_110000000000000000000000
Q = 125 / 6 = 20 = 000000000000000000010100
REM = 5 = 000000000000000000000101

根据Divisor的值, 可得选择常数:
m[-1] 	= -19 	= 110_1101
m[0] 	= -6 	= 111_1001
m[1] 	= 6		= 000_0110
m[2] 	= 19	= 001_0011

D = 000_11000000000000000000000000
2D = 001_10000000000000000000000000
-D = 111_01000000000000000000000000
-2D = 110_10000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[3] = 1_11100000000000000000000000 < 0
q[final] = q[3]
q_pos = 0101_01
q_neg = 0000_00
q_calculated_pre = q_pos - q_neg = 010101
q_calculated = q_calculated_pre - (w[final] < 0) = 010100
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
(111000000000000000000000 + 110000000000000000000000) >> 21 = 
101000000000000000000000 >> 21 = 
000000000000000000000101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00111110100000000000000000
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 10
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_11111010000000000000000000 + 
111_01000000000000000000000000 = 
000_00111010000000000000000000 -> 
w[1] = 0_00111010000000000000000000
4 * w[1] = 000_11101000000000000000000000
(4 * w[1])_trunc_3_4 = 000_1110, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 1010
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_11101000000000000000000000 + 
111_01000000000000000000000000 = 
000_00101000000000000000000000 -> 
w[2] = 0_00101000000000000000000000
4 * w[2] = 000_10100000000000000000000000
(4 * w[2])_trunc_3_4 = 000_1010, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0101_01
q_neg = 0000_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_10100000000000000000000000 + 
111_01000000000000000000000000 = 
111_11100000000000000000000000 -> 
w[3] = 1_11100000000000000000000000
4 * w[3] = 111_10000000000000000000000000
(4 * w[3])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0101_0100
q_neg = 0000_0001


// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 000000000101011110000000 = 22400
D[24-1:0] = 000000000000000000001100 = 12
Q[24-1:0] = X / D = 1866 = 000000000000011101001010
REM[24-1:0] = 22400 - 12 * 1866 = 8 = 000000000000000000001000
按照小数除法的方式, 将X和D规格化:
CLZ_X = 9
CLZ_D = 20
CLZ_DIFF = CLZ_D - CLZ_X = 11
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 7
CLZ_DIFF为奇数 -> 将Dividend规格化到区间"[1/4, 1/2)"上
Dividend[25-1:0] 	= 0_010101111000000000000000
Divisor[25-1:0] 	= 0_110000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -19 	= 110_1101
m[0] 	= -6 	= 111_1001
m[1] 	= 6		= 000_0110
m[2] 	= 19	= 001_0011

+ D = 000_11000000000000000000000000
+2D = 001_10000000000000000000000000
- D = 111_01000000000000000000000000
-2D = 110_10000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[7] = 1_11000000000000000000000000 < 0
q[final] = q[7]
q_pos = 0010_0001_0100_00
q_neg = 0000_0100_0001_01
q_calculated_pre = q_pos - q_neg = 011101001011
q_calculated = q_calculated_pre - (w[final] < 0) = 011101001010
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
(110000000000000000000000 + 110000000000000000000000) >> 20 = 
100000000000000000000000 >> 20 = 
000000000000000000001000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00010101111000000000000000
4 * w[0] = 000_01010111100000000000000000
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_0101, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_01010111100000000000000000 + 
000_00000000000000000000000000 = 
000_01010111100000000000000000 -> 
w[1] = 0_01010111100000000000000000
4 * w[1] = 001_01011110000000000000000000
(4 * w[1])_trunc_3_4 = 001_0101, "belongs to [m[2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
001_01011110000000000000000000 + 
110_10000000000000000000000000 = 
111_11011110000000000000000000 -> 
w[2] = 1_11011110000000000000000000
4 * w[2] = 111_01111000000000000000000000
(4 * w[2])_trunc_3_4 = 111_0111, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0010_00
q_neg = 0000_01

ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_01111000000000000000000000 + 
000_11000000000000000000000000 = 
000_00111000000000000000000000 -> 
w[3] = 0_00111000000000000000000000
4 * w[3] = 000_11100000000000000000000000
(4 * w[3])_trunc_3_4 = 000_1110, "belongs to [m[1], m[2])" -> q[4] = +1
q_pos = 0010_0001
q_neg = 0000_0100

ITER[3]:
4 * w[3] + (-q[4] * D) = 
000_11100000000000000000000000 + 
111_01000000000000000000000000 = 
000_00100000000000000000000000 -> 
w[4] = 0_00100000000000000000000000
4 * w[4] = 000_10000000000000000000000000
(4 * w[4])_trunc_3_4 = 000_1000, "belongs to [m[1], m[2])" -> q[5] = +1
q_pos = 0010_0001_01
q_neg = 0000_0100_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
000_10000000000000000000000000 + 
111_01000000000000000000000000 = 
111_11000000000000000000000000 -> 
w[5] = 1_11000000000000000000000000
4 * w[5] = 111_00000000000000000000000000
(4 * w[5])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0010_0001_0100
q_neg = 0000_0100_0001

// 从现在开始进入循环...
ITER[5]:
4 * w[5] + (-q[6] * D) = 
111_00000000000000000000000000 + 
000_11000000000000000000000000 = 
111_11000000000000000000000000 -> 
w[6] = 1_11000000000000000000000000
4 * w[6] = 111_00000000000000000000000000
(4 * w[6])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0010_0001_0100_00
q_neg = 0000_0100_0001_01

ITER[6]:
4 * w[6] + (-q[7] * D) = 
111_00000000000000000000000000 + 
000_11000000000000000000000000 = 
111_11000000000000000000000000 -> 
w[7] = 1_11000000000000000000000000
4 * w[7] = 111_00000000000000000000000000
(4 * w[7])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[8] = -1
q_pos = 0010_0001_0100_0000
q_neg = 0000_0100_0001_0101

// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 000000000101011110000111 = 22407
D[24-1:0] = 000000000000000010111001 = 185
Q[24-1:0] = X / D = 121 = 000000000000000001111001
REM[24-1:0] = 22407 - 185 * 121 = 22 = 000000000000000000010110
按照小数除法的方式, 将X和D规格化:
CLZ_X = 9
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 7
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 5
CLZ_DIFF为奇数 -> 将Dividend规格化到区间"[1/4, 1/2)"上
Dividend[25-1:0] 	= 0_010101111000011100000000
Divisor[25-1:0] 	= 0_101110010000000000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -17 	= 110_1111
m[0] 	= -6 	= 111_1001
m[1] 	= 6		= 000_0110
m[2] 	= 17	= 001_0001

D = 000_10111001000000000000000000
2D = 001_01110010000000000000000000
-D = 111_01000111000000000000000000
-2D = 110_10001110000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[5] = 0_00010110000000000000000000 > 0
q[final] = q[5]:
q_pos = 0010_0000_01
q_neg = 0000_0010_00
q_calculated_pre = q_pos - q_neg = 01111001
q_calculated = q_calculated_pre - (w[final]< 0) = 01111001 = 01111001
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
000101100000000000000000 >> 16 = 
000000000000000000010110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00010101111000011100000000
4 * w[0] = 000_01010111100001110000000000
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_0101, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_01010111100001110000000000 + 
000_00000000000000000000000000 = 
000_01010111100001110000000000 -> 
w[1] = 0_01010111100001110000000000
4 * w[1] = 001_01011110000111000000000000
(4 * w[1])_trunc_3_4 = 001_0101, "belongs to [m[2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
001_01011110000111000000000000 + 
110_10001110000000000000000000 = 
111_11101100000111000000000000 -> 
w[2] = 1_11101100000111000000000000
4 * w[2] = 111_10110000011100000000000000
(4 * w[2])_trunc_3_4 = 111_1011, "belongs to [m[0], m[1])" -> q[3] = 0
q_pos = 0010_00
q_neg = 0000_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_10110000011100000000000000 + 
000_00000000000000000000000000 = 
111_10110000011100000000000000 -> 
w[3] = 1_10110000011100000000000000
4 * w[3] = 110_11000001110000000000000000
(4 * w[3])_trunc_3_4 = 110_1100, "belongs to [-Inf, m[-1])" -> q[4] = -2
q_pos = 0010_0000
q_neg = 0000_0010

ITER[3]:
4 * w[3] + (-q[4] * D) = 
110_11000001110000000000000000 + 
001_01110010000000000000000000 = 
000_00110011110000000000000000 -> 
w[4] = 0_00110011110000000000000000
4 * w[4] = 000_11001111000000000000000000
(4 * w[4])_trunc_3_4 = 000_1100, "belongs to [m[1], m[2])" -> q[5] = +1
q_pos = 0010_0000_01
q_neg = 0000_0010_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
000_11001111000000000000000000 + 
111_01000111000000000000000000 = 
000_00010110000000000000000000 -> 
w[5] = 0_00010110000000000000000000
4 * w[5] = 000_01011000000000000000000000
(4 * w[5])_trunc_3_4 = 000_0101, "belongs to [m[0], m[1])" -> q[6] = 0
q_pos = 0010_0000_0100
q_neg = 0000_0010_0000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 000000111101011110000011 = 251779
D[24-1:0] = 000000000000000110101011 = 427
Q[24-1:0] = X / D = 589 = 000000000000001001001101
REM[24-1:0] = 251779 - 427 * 589 = 276 = 000000000000000100010100
按照小数除法的方式, 将X和D规格化:
CLZ_X = 6
CLZ_D = 15
CLZ_DIFF = CLZ_D - CLZ_X = 9
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 6
CLZ_DIFF为奇数 -> 将Dividend规格化到区间"[1/4, 1/2)"上
Dividend[25-1:0] 	= 0_011110101111000001100000
Divisor[25-1:0] 	= 0_110101011000000000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -20 	= 110_1100
m[0] 	= -6 	= 111_1001
m[1] 	= 6		= 000_0110
m[2] 	= 20	= 001_0100

D = 000_11010101100000000000000000
2D = 001_10101011000000000000000000
-D = 111_00101010100000000000000000
-2D = 110_01010101000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[6] = 1_10110100100000000000000000 < 0
q[final] = q[6]:
q_pos = 0100_0101_0010
q_neg = 0010_0000_0100
q_calculated_pre = q_pos - q_neg = 001001001110
q_calculated = q_calculated_pre - (w[final] < 0) = 001001001110 = 001001001101
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
(101101001000000000000000 + 110101011000000000000000) >> 15 = 
100010100000000000000000 >> 15
000000000000000100010100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][27-1:0] = Dividend / 4 = 0_00011110101111000001100000
4 * w[0] = 000_01111010111100000110000000
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_0111, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_01111010111100000110000000 + 
111_00101010100000000000000000 = 
111_10100101011100000110000000 -> 
w[1] = 1_10100101011100000110000000
4 * w[1] = 110_10010101110000011000000000
(4 * w[1])_trunc_3_4 = 110_1001, "belongs to [-Inf, m[-1])" -> q[2] = -2
q_pos = 0100
q_neg = 0010

ITER[1]:
4 * w[1] + (-q[2] * D) = 
110_10010101110000011000000000 + 
001_10101011000000000000000000 = 
000_01000000110000011000000000 -> 
w[2] = 0_01000000110000011000000000
4 * w[2] = 001_00000011000001100000000000
(4 * w[2])_trunc_3_4 = 001_0000, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0100_01
q_neg = 0010_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
001_00000011000001100000000000 + 
111_00101010100000000000000000 = 
000_00101101100001100000000000 -> 
w[3] = 0_00101101100001100000000000
4 * w[3] = 000_10110110000110000000000000
(4 * w[3])_trunc_3_4 = 000_1011, "belongs to [m[1], m[2])" -> q[4] = +1
q_pos = 0100_0101
q_neg = 0010_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
000_10110110000110000000000000 + 
111_00101010100000000000000000 = 
111_11100000100110000000000000 -> 
w[4] = 1_11100000100110000000000000
4 * w[4] = 111_10000010011000000000000000
(4 * w[4])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[5] = -1
q_pos = 0100_0101_00
q_neg = 0010_0000_01

ITER[4]:
4 * w[4] + (-q[5] * D) = 
111_10000010011000000000000000 + 
000_11010101100000000000000000 = 
000_01010111111000000000000000 -> 
w[5] = 0_01010111111000000000000000
4 * w[5] = 001_01011111100000000000000000
(4 * w[5])_trunc_3_4 = 001_0101, "belongs to [m[2], +Inf)" -> q[6] = +2
q_pos = 0100_0101_0010
q_neg = 0010_0000_0100

ITER[5]:
4 * w[5] + (-q[6] * D) = 
001_01011111100000000000000000 + 
110_01010101000000000000000000 = 
111_10110100100000000000000000 -> 
w[6] = 1_10110100100000000000000000
4 * w[6] = 110_11010010000000000000000000
(4 * w[6])_trunc_3_4 = 110_1101, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0100_0101_0010_00
q_neg = 0010_0000_0100_01

// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 010011110101011110000111 = 5199751
D[24-1:0] = 000000000000000001110100 = 116
Q[24-1:0] = X / D = 44825 = 000000001010111100011001
REM[24-1:0] = 5199751 - 116 * 44825 = 51 = 000000000000000000110011
按照小数除法的方式, 将X和D规格化:
CLZ_X = 1
CLZ_D = 17
CLZ_DIFF = CLZ_D - CLZ_X = 16
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 9
Dividend[25-1:0] 	= 0_100111101010111100001110
Divisor[25-1:0] 	= 0_111010000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -22 	= 110_1010
m[0] 	= -8 	= 111_1000
m[1] 	= 8		= 000_1000
m[2] 	= 22	= 001_0110

D = 000_11101000000000000000000000
2D = 001_11010000000000000000000000
-D = 111_00011000000000000000000000
-2D = 110_00110000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[9] = 0_01100110000000000000000000 > 0
q[final] = q[9]:
q_pos = 0100_0000_0000_1000_01
q_neg = 0001_0100_0100_0010_00
q_calculated_pre = q_pos - q_neg = 1010111100011001
q_calculated = q_calculated_pre - (w[final] < 0) = 1010111100011001
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
011001100000000000000000 >> 17 = 
000000000000000000110011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00100111101010111100001110
4 * w[0] = 000_10011110101011110000111000
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_1001, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_10011110101011110000111000 + 
111_00011000000000000000000000 = 
111_10110110101011110000111000 -> 
w[1] = 1_10110110101011110000111000
4 * w[1] = 110_11011010101111000011100000
(4 * w[1])_trunc_3_4 = 110_1101, "belongs to [m[-1], m[0])" -> q[2] = -1
q_pos = 0100
q_neg = 0001

ITER[1]:
4 * w[1] + (-q[2] * D) = 
110_11011010101111000011100000 + 
000_11101000000000000000000000 = 
111_11000010101111000011100000 -> 
w[2] = 1_11000010101111000011100000
4 * w[2] = 111_00001010111100001110000000
(4 * w[2])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0100_00
q_neg = 0001_01

ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_00001010111100001110000000 + 
000_11101000000000000000000000 = 
111_11110010111100001110000000 -> 
w[3] = 1_11110010111100001110000000
4 * w[3] = 111_11001011110000111000000000
(4 * w[3])_trunc_3_4 = 111_1100, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0100_0000
q_neg = 0001_0100

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_11001011110000111000000000 + 
000_00000000000000000000000000 = 
111_11001011110000111000000000 -> 
w[4] = 1_11001011110000111000000000
4 * w[4] = 111_00101111000011100000000000
(4 * w[4])_trunc_3_4 = 111_0010, "belongs to [m[-1], m[0])" -> q[5] = -1
q_pos = 0100_0000_00
q_neg = 0001_0100_01

ITER[4]:
4 * w[4] + (-q[5] * D) = 
111_00101111000011100000000000 + 
000_11101000000000000000000000 = 
000_00010111000011100000000000 -> 
w[5] = 0_00010111000011100000000000
4 * w[5] = 000_01011100001110000000000000
(4 * w[5])_trunc_3_4 = 000_0101, "belongs to [m[0], m[1])" -> q[6] = 0
q_pos = 0100_0000_0000
q_neg = 0001_0100_0100

ITER[5]:
4 * w[5] + (-q[6] * D) = 
000_01011100001110000000000000 + 
000_00000000000000000000000000 = 
000_01011100001110000000000000 -> 
w[6] = 0_01011100001110000000000000
4 * w[6] = 001_01110000111000000000000000
(4 * w[6])_trunc_3_4 = 001_0111, "belongs to [m[2], +Inf)" -> q[7] = +2
q_pos = 0100_0000_0000_10
q_neg = 0001_0100_0100_00

ITER[6]:
4 * w[6] + (-q[7] * D) = 
001_01110000111000000000000000 + 
110_00110000000000000000000000 = 
111_10100000111000000000000000 -> 
w[7] = 1_10100000111000000000000000
4 * w[7] = 110_10000011100000000000000000
(4 * w[7])_trunc_3_4 = 110_1000, "belongs to [-Inf, m[-1])" -> q[8] = -2
q_pos = 0100_0000_0000_1000
q_neg = 0001_0100_0100_0010

ITER[7]:
4 * w[7] + (-q[8] * D) = 
110_10000011100000000000000000 + 
001_11010000000000000000000000 = 
000_01010011100000000000000000 -> 
w[8] = 0_01010011100000000000000000
4 * w[8] = 001_01001110000000000000000000
(4 * w[8])_trunc_3_4 = 001_0100, "belongs to [m[1], m[2])" -> q[9] = +1
q_pos = 0100_0000_0000_1000_01
q_neg = 0001_0100_0100_0010_00

ITER[8]:
4 * w[8] + (-q[9] * D) = 
001_01001110000000000000000000 + 
111_00011000000000000000000000 = 
000_01100110000000000000000000 -> 
w[9] = 0_01100110000000000000000000
4 * w[9] = 001_10011000000000000000000000
(4 * w[9])_trunc_3_4 = 001_1001, "belongs to [m[2], +Inf)" -> q[10] = +2
q_pos = 0100_0000_0000_1000_0110
q_neg = 0001_0100_0100_0010_0000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[24-1:0] = 010010011001111001100111 = 4824679
D[24-1:0] = 000000000000000011000101 = 197
Q[24-1:0] = X / D = 24490 = 000000000101111110101010
REM[24-1:0] = 4824679 - 197 * 24490 = 149 = 000000000000000010010101
按照小数除法的方式, 将X和D规格化:
CLZ_X = 1
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 15
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / 2) = 9
CLZ_DIFF为奇数 -> 将Dividend规格化到区间"[1/4, 1/2)"上
Dividend[25-1:0] 	= 0_010010011001111001100111
Divisor[25-1:0] 	= 0_110001010000000000000000
根据Divisor的值, 可得选择常数:
m[-1] 	= -19 	= 110_1101
m[0] 	= -6 	= 111_1001
m[1] 	= 6		= 000_0110
m[2] 	= 19	= 001_0011

D = 000_11000101000000000000000000
2D = 001_10001010000000000000000000
-D = 111_00111011000000000000000000
-2D = 110_01110110000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
w[final] = w[9] = 1_11010000000000000000000000 < 0
q[final] = q[9]:
q_pos = 0001_1000_0000_0000_00
q_neg = 0000_0000_0001_0101_01
q_calculated_pre = q_pos - q_neg = 0101111110101011
q_calculated = q_calculated_pre - (w[final] < 0) = 0101111110101011 = 0101111110101010
remainder = (w[final][2 +: 24] + ((w[final] < 0) ? Divisor : 24'b0)) >> CLZ_D = 
(110100000000000000000000 + 110001010000000000000000) >> 16 = 
100101010000000000000000 >> 16 = 
000000000000000010010101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][27-1:0] = Dividend / 4 = 0_00010010011001111001100111
4 * w[0] = 000_01001001100111100110011100
q[0] = 0
(4 * w[0])_trunc_3_4 = 000_0100, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_01001001100111100110011100 + 
000_00000000000000000000000000 = 
000_01001001100111100110011100 -> 
w[1] = 0_01001001100111100110011100
4 * w[1] = 001_00100110011110011001110000
(4 * w[1])_trunc_3_4 = 001_0010, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
001_00100110011110011001110000 + 
111_00111011000000000000000000 = 
000_01100001011110011001110000 -> 
w[2] = 0_01100001011110011001110000
4 * w[2] = 001_10000101111001100111000000
(4 * w[2])_trunc_3_4 = 001_1000, "belongs to [m[2], +Inf)" -> q[3] = +2
q_pos = 0001_10
q_neg = 0000_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
001_10000101111001100111000000 + 
110_01110110000000000000000000 = 
111_11111011111001100111000000 -> 
w[3] = 1_11111011111001100111000000
4 * w[3] = 111_11101111100110011100000000
(4 * w[3])_trunc_3_4 = 111_1110, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0001_1000
q_neg = 0000_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_11101111100110011100000000 + 
000_00000000000000000000000000 = 
111_11101111100110011100000000 -> 
w[4] = 1_11101111100110011100000000
4 * w[4] = 111_10111110011001110000000000
(4 * w[4])_trunc_3_4 = 111_1011, "belongs to [m[0], m[1])" -> q[5] = 0
q_pos = 0001_1000_00
q_neg = 0000_0000_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
111_10111110011001110000000000 + 
000_00000000000000000000000000 = 
111_10111110011001110000000000 -> 
w[5] = 1_10111110011001110000000000
4 * w[5] = 110_11111001100111000000000000
(4 * w[5])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0001_1000_0000
q_neg = 0000_0000_0001

ITER[5]:
4 * w[5] + (-q[6] * D) = 
110_11111001100111000000000000 + 
000_11000101000000000000000000 = 
111_10111110100111000000000000 -> 
w[6] = 1_10111110100111000000000000
4 * w[6] = 110_11111010011100000000000000
(4 * w[6])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0001_1000_0000_00
q_neg = 0000_0000_0001_01

ITER[6]:
4 * w[6] + (-q[7] * D) = 
110_11111010011100000000000000 + 
000_11000101000000000000000000 = 
111_10111111011100000000000000 -> 
w[7] = 1_10111111011100000000000000
4 * w[7] = 110_11111101110000000000000000
(4 * w[7])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[8] = -1
q_pos = 0001_1000_0000_0000
q_neg = 0000_0000_0001_0101

ITER[7]:
4 * w[7] + (-q[8] * D) = 
110_11111101110000000000000000 + 
000_11000101000000000000000000 = 
111_11000010110000000000000000 -> 
w[8] = 1_11000010110000000000000000
4 * w[8] = 111_00001011000000000000000000
(4 * w[8])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[9] = -1
q_pos = 0001_1000_0000_0000_00
q_neg = 0000_0000_0001_0101_01

ITER[8]:
4 * w[8] + (-q[9] * D) = 
111_00001011000000000000000000 + 
000_11000101000000000000000000 = 
111_11010000000000000000000000 -> 
w[9] = 1_11010000000000000000000000
4 * w[9] = 111_01000000000000000000000000
(4 * w[9])_trunc_3_4 = 111_0100, "belongs to [m[-1], m[0])" -> q[10] = -1
q_pos = 0001_1000_0000_0000_0000
q_neg = 0000_0000_0001_0101_0101






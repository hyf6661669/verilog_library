测试MultiCycle-Path形式实现的Radix-4 SRT除法.
对于"CLZ_D = WIDTH - 1"的情况(即divisor = {(WIDTH - 1){1'b0}, 1'b1})，不通过迭代的方式得到最终的结果，而是将其视为特殊情况，和"divisor_is_zero"信号一起通过Mux来生成输出信号.


// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 24;
ITN = InTerNal
ITN_W = 1 + (2 * WIDTH) = 49;
0_000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 100010101001010010010100 = 9082004
D[WIDTH-1:0] = 100000000000000000000011 = 8388611
Q[WIDTH-1:0] = X / D = 1 = 000000000000000000000001
REM[WIDTH-1:0] = 9082004 - 1 * 8388611 = 693393 = 000010101001010010010001

CLZ_X = 0
CLZ_D = 0
CLZ_DIFF = CLZ_D - CLZ_X = 0
Normalized_D = 100000000000000000000011
根据D的值, 可得选择常数:
m[-1] = -18
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

+ D = 0_100000000000000000000011
+2D = 1_000000000000000000000110
- D = 1_011111111111111111111101
-2D = 0_111111111111111111111010

l_shift_num = CLZ_D = 0
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_000000000000000000000000100010101001010010010100 << 0 = 
0_000000000000000000000000100010101001010010010100

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:WIDTH] = 0_000000000000000000000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
100010101001010010010100

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_000000000000000000000010 + 
0_000000000000000000000000 = 
0_000000000000000000000010
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
001010100101001001010000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_000000000000000000001000 + 
0_000000000000000000000000 = 
0_000000000000000000001000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
101010010100100101000000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_000000000000000000100010 + 
0_000000000000000000000000 = 
0_000000000000000000100010
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
101001010010010100000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_000000000000000010001010 + 
0_000000000000000000000000 = 
0_000000000000000010001010
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
100101001001010000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_000000000000001000101010 + 
0_000000000000000000000000 = 
0_000000000000001000101010
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
010100100101000000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_000000000000100010101001 + 
0_000000000000000000000000 = 
0_000000000000100010101001
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
010010010100000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_000000000010001010100101 + 
0_000000000000000000000000 = 
0_000000000010001010100101
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
001001010000000000000000

ITER[7]:
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_000000001000101010010100 + 
0_000000000000000000000000 = 
0_000000001000101010010100
(4 * w[8])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
100101000000000000000000

ITER[8]:
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_000000100010101001010010 + 
0_000000000000000000000000 = 
0_000000100010101001010010
(4 * w[9])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
010100000000000000000000

ITER[9]:
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_000010001010100101001001 + 
0_000000000000000000000000 = 
0_000010001010100101001001
(4 * w[10])_trunc_3_4 = 000_0010, "belongs to [m[0], m[+1])" -> q[11] = 0
q_pos = 0000_0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
010000000000000000000000

ITER[10]:
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
0_001000101010010100100101 + 
0_000000000000000000000000 = 
0_001000101010010100100101
(4 * w[11])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[12] = +1
q_pos = 0000_0000_0000_0000_0000_0001
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[12] = {w[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[12] * D = 
0_100010101001010010010100 + 
1_011111111111111111111101 = 
0_000010101001010010010001 >= 0

rem = (w[12])_reduced >> CLZ_D = 
000010101001010010010001 >> 0
000010101001010010010001

q_final = corr(q_pos - q_neg) = 000000000000000000000001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 24;
ITN = InTerNal
ITN_W = 1 + (2 * WIDTH) = 49;
0000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 100010101001010010010100 = 9082004
D[WIDTH-1:0] = 000000000000000000000011 = 3
Q[WIDTH-1:0] = X / D = 3027334 = 001011100011000110000110
REM[WIDTH-1:0] = 9082004 - 3 * 3027334 = 2 = 000000000000000000000010

CLZ_X = 0
CLZ_D = 22
CLZ_DIFF = CLZ_D - CLZ_X = 22
Normalized_D = 110000000000000000000000
根据D的值, 可得选择常数:
m[-1] = -18
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

+ D = 0_110000000000000000000000
+2D = 1_100000000000000000000000
- D = 1_010000000000000000000000
-2D = 0_100000000000000000000000

l_shift_num = CLZ_D = 22
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_000000000000000000000000100010101001010010010100 << 22 = 
0_001000101010010100100101000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:WIDTH] = 0_001000101010010100100101
(4 * w[0])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
000000000000000000000000

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_100010101001010010010100 + 
1_010000000000000000000000 = 
1_110010101001010010010100
(4 * w[1])_trunc_3_4 = 111_0010, "belongs to [m[-1], m[0])" -> q[2] = -1
q_pos = 0100
q_neg = 0001
temp_dividend[1] = temp_dividend[0] << 2 = 
000000000000000000000000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
1_001010100101001001010000 + 
0_110000000000000000000000 = 
1_111010100101001001010000
(4 * w[2])_trunc_3_4 = 111_1010, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0100_00
q_neg = 0001_00
temp_dividend[2] = temp_dividend[1] << 2 = 
000000000000000000000000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
1_101010010100100101000000 + 
0_000000000000000000000000 = 
1_101010010100100101000000
(4 * w[3])_trunc_3_4 = 110_1010, "belongs to [-Inf, m[-1])" -> q[4] = -2
q_pos = 0100_0000
q_neg = 0001_0010
temp_dividend[3] = temp_dividend[2] << 2 = 
000000000000000000000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_101001010010010100000000 + 
1_100000000000000000000000 = 
0_001001010010010100000000
(4 * w[4])_trunc_3_4 = 000_1001, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0100_0000_01
q_neg = 0001_0010_00
temp_dividend[4] = temp_dividend[3] << 2 = 
000000000000000000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_100101001001010000000000 + 
1_010000000000000000000000 = 
1_110101001001010000000000
(4 * w[5])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0100_0000_0100
q_neg = 0001_0010_0001
temp_dividend[5] = temp_dividend[4] << 2 = 
000000000000000000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
1_010100100101000000000000 + 
0_110000000000000000000000 = 
0_000100100101000000000000
(4 * w[6])_trunc_3_4 = 000_0100, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0100_0000_0100_00
q_neg = 0001_0010_0001_00
temp_dividend[6] = temp_dividend[5] << 2 = 
000000000000000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_010010010100000000000000 + 
0_000000000000000000000000 = 
0_010010010100000000000000
(4 * w[7])_trunc_3_4 = 001_0010, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0100_0000_0100_0010
q_neg = 0001_0010_0001_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
000000000000000000000000

ITER[7]:
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
1_001001010000000000000000 + 
0_100000000000000000000000 = 
1_101001010000000000000000
(4 * w[8])_trunc_3_4 = 110_1001, "belongs to [-Inf, m[-1])" -> q[9] = -2
q_pos = 0100_0000_0100_0010_00
q_neg = 0001_0010_0001_0000_10
temp_dividend[8] = temp_dividend[7] << 2 = 
000000000000000000000000

ITER[8]:
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_100101000000000000000000 + 
1_100000000000000000000000 = 
0_000101000000000000000000
(4 * w[9])_trunc_3_4 = 000_0101, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0100_0000_0100_0010_0000
q_neg = 0001_0010_0001_0000_1000
temp_dividend[9] = temp_dividend[8] << 2 = 
000000000000000000000000

ITER[9]:
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_010100000000000000000000 + 
0_000000000000000000000000 = 
0_010100000000000000000000
(4 * w[10])_trunc_3_4 = 001_0100, "belongs to [m[+2], +Inf)" -> q[11] = +2
q_pos = 0100_0000_0100_0010_0000_10
q_neg = 0001_0010_0001_0000_1000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
000000000000000000000000

ITER[10]:
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
1_010000000000000000000000 + 
0_100000000000000000000000 = 
1_110000000000000000000000
(4 * w[11])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[12] = -1
q_pos = 0100_0000_0100_0010_0000_1000
q_neg = 0001_0010_0001_0000_1000_0001
temp_dividend[11] = temp_dividend[10] << 2 = 
000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[12] = {w[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[12] * D = 
1_000000000000000000000000 + 
0_110000000000000000000000 = 
1_110000000000000000000000 < 0

rem = (w[12] + D)_reduced >> CLZ_D = 
(110000000000000000000000 + 110000000000000000000000) >> 22 = 
100000000000000000000000 >> 22 = 
000000000000000000000010

q_final = corr(q_pos - q_neg) = 001011100011000110000110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 100010101001010010010100 = 9082004
D[WIDTH-1:0] = 000100110011001110001001 = 1258377
Q[WIDTH-1:0] = X / D = 7 = 000000000000000000000111
REM[WIDTH-1:0] = 9082004 - 1258377 * 7 = 273365 = 000001000010101111010101

CLZ_X = 0
CLZ_D = 3
CLZ_DIFF = CLZ_D - CLZ_X = 3
Normalized_D = 100110011001110001001000
根据D的值, 可得选择常数:
m[-1] = -14
m[ 0] = - 4
m[+1] = + 4
m[+2] = +14

+ D = 0_100110011001110001001000
+2D = 1_001100110011100010010000
- D = 1_011001100110001110111000
-2D = 0_110011001100011101110000

l_shift_num = CLZ_D = 3
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_000000000000000000000000100010101001010010010100 << 3 = 
0_000000000000000000000100010101001010010010100000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:WIDTH] = 0_000000000000000000000100
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
010101001010010010100000

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_000000000000000000010001 + 
0_000000000000000000000000 = 
0_000000000000000000010001
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
010100101001001010000000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_000000000000000001000101 + 
0_000000000000000000000000 = 
0_000000000000000001000101
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
010010100100101000000000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_000000000000000100010101 + 
0_000000000000000000000000 = 
0_000000000000000100010101
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
001010010010100000000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_000000000000010001010100 + 
0_000000000000000000000000 = 
0_000000000000010001010100
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
101001001010000000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_000000000001000101010010 + 
0_000000000000000000000000 = 
0_000000000001000101010010
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
100100101000000000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_000000000100010101001010 + 
0_000000000000000000000000 = 
0_000000000100010101001010
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
010010100000000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_000000010001010100101001 + 
0_000000000000000000000000 = 
0_000000010001010100101001
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
001010000000000000000000

ITER[7]:
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_000001000101010010100100 + 
0_000000000000000000000000 = 
0_000001000101010010100100
(4 * w[8])_trunc_3_4 = 000_0001, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
101000000000000000000000

ITER[8]:
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_000100010101001010010010 + 
0_000000000000000000000000 = 
0_000100010101001010010010
(4 * w[9])_trunc_3_4 = 000_0100, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
100000000000000000000000

ITER[9]:
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_010001010100101001001010 + 
0_000000000000000000000000 = 
0_010001010100101001001010
(4 * w[10])_trunc_3_4 = 001_0001, "belongs to [m[0], m[+1])" -> q[11] = +2
q_pos = 0000_0000_0000_0000_0000_10
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
000000000000000000000000

ITER[10]:
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
1_000101010010100100101000 + 
0_110011001100011101110000 = 
1_111000011111000010011000
(4 * w[11])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[12] = 0
q_pos = 0000_0000_0000_0000_0000_1000
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[12] = {w[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[12] * D = 
1_100001111100001001100000 + 
0_000000000000000000000000 = 
1_100001111100001001100000 < 0

rem = (w[12] + D)_reduced >> CLZ_D = 
(100001111100001001100000 + 100110011001110001001000) >> 3
001000010101111010101000 >> 3 = 
000001000010101111010101

q_final = corr(q_pos - q_neg) = 000000000000000000000111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000000000000000000101000 = 40
D[WIDTH-1:0] = 000000000111101110001110 = 31630
Q[WIDTH-1:0] = X / D = 0 = 000000000000000000000000
REM[WIDTH-1:0] = 40 - 31630 * 0 = 40 = 000000000000000000101000

CLZ_X = 18
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = -9
Normalized_D = 111101110001110000000000
根据D的值, 可得选择常数:
m[-1] = -23
m[ 0] = - 8
m[+1] = + 8
m[+2] = +23

+ D = 0_111101110001110000000000
+2D = 1_111011100011100000000000
- D = 1_000010001110010000000000
-2D = 0_000100011100100000000000

l_shift_num = CLZ_D = 9
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_000000000000000000000000000000000000000000101000 << 9 = 
0_000000000000000000000000000000000101000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:WIDTH] = 0_000000000000000000000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
000000000101000000000000

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_000000000000000000000000 + 
0_000000000000000000000000 = 
0_000000000000000000000000
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
000000010100000000000000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_000000000000000000000000 + 
0_000000000000000000000000 = 
0_000000000000000000000000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
000001010000000000000000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_000000000000000000000000 + 
0_000000000000000000000000 = 
0_000000000000000000000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
000101000000000000000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_000000000000000000000000 + 
0_000000000000000000000000 = 
0_000000000000000000000000
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
010100000000000000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_000000000000000000000001 + 
0_000000000000000000000000 = 
0_000000000000000000000001
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
010000000000000000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_000000000000000000000101 + 
0_000000000000000000000000 = 
0_000000000000000000000101
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
000000000000000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_000000000000000000010100 + 
0_000000000000000000000000 = 
0_000000000000000000010100
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
000000000000000000000000

ITER[7]:
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_000000000000000001010000 + 
0_000000000000000000000000 = 
0_000000000000000001010000
(4 * w[8])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
000000000000000000000000

ITER[8]:
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_000000000000000101000000 + 
0_000000000000000000000000 = 
0_000000000000000101000000
(4 * w[9])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
000000000000000000000000

ITER[9]:
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_000000000000010100000000 + 
0_000000000000000000000000 = 
0_000000000000010100000000
(4 * w[10])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[11] = 0
q_pos = 0000_0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
000000000000000000000000

ITER[10]:
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
0_000000000001010000000000 + 
0_000000000000000000000000 = 
0_000000000001010000000000
(4 * w[11])_trunc_3_4 = 000_0000, "belongs to [m[-1], m[0])" -> q[12] = 0
q_pos = 0000_0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[12] = {w[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[12] * D = 
0_000000000101000000000000 + 
0_000000000000000000000000 = 
0_000000000101000000000000 >= 0

rem = (w[12])_reduced >> CLZ_D = 
000000000101000000000000 >> 9 = 
000000000000000000101000

q_final = corr(q_pos - q_neg) = 000000000000000000000000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------








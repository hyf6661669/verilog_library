// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 11111101000011100111001000110000 = 4245582384
D[WIDTH-1:0] = 11100000000101000000000010000000 = 3759407232
Q[WIDTH-1:0] = X / D = 1 = 00000000000000000000000000000001
REM[WIDTH-1:0] = 4245582384 - 3759407232 * 1 = 486175152 = 00011100111110100111000110110000

CLZ_X = 0
CLZ_D = 0
CLZ_DIFF = CLZ_D - CLZ_X = 0
r_shift_num = CLZ_DIFF[0] = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(2 / 2) = 1;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11111101000011100111001000110000
Divisor[WIDTH-1:0] 		= 11100000000101000000000010000000

+ D = 0_11100000000101000000000010000000000
+2D = 1_11000000001010000000000100000000000
- D = 1_00011111111010111111111110000000000
-2D = 0_00111111110101111111111100000000000
~ D = 1_00011111111010111111111101111111111
~2D = 0_00111111110101111111111011111111111

根据D的值, 可得选择常数:
m[-1] = -22
m[ 0] = - 8
m[+1] = + 8 = 00_1000
m[+2] = +22 = 01_0110

// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0] = 0_00111111010000111001110010001100000

(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

csa_3_2_x1 = 0_11111101000011100111001000110000000

w[1] = 4 * w[0] - q[1] * D = 
0_11111101000011100111001000110000000 + 
1_00011111111010111111111110000000000 = 
0_00011100111110100111000110110000000

w[1]_reduced >> CLZ_D = 
00011100111110100111000110110000

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 11111101000011100111001000110000 = 4245582384
D[WIDTH-1:0] = 01110000000010100000000001000000 = 1879703616
Q[WIDTH-1:0] = X / D = 2 = 00000000000000000000000000000010
REM[WIDTH-1:0] = 4245582384 - 1879703616 * 2 = 486175152 = 00011100111110100111000110110000

CLZ_X = 0
CLZ_D = 1
CLZ_DIFF = CLZ_D - CLZ_X = 1
r_shift_num = CLZ_DIFF[0] = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(3 / 2) = 2;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11111101000011100111001000110000
Divisor[WIDTH-1:0] 		= 11100000000101000000000010000000

+ D = 0_11100000000101000000000010000000000
+2D = 1_11000000001010000000000100000000000
- D = 1_00011111111010111111111110000000000
-2D = 0_00111111110101111111111100000000000

根据D的值, 可得选择常数:
m[-1] = -22
m[ 0] = - 8
m[+1] = + 8
m[+2] = +22

// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0] = 0_00011111101000011100111001000110000
(4 * w[0])_trunc_3_4 = 000_0111, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

w[1] = 4 * w[0] - q[1] * D = 
0_01111110100001110011100100011000000 + 
0_00000000000000000000000000000000000 = 
0_01111110100001110011100100011000000
(4 * w[1])_trunc_3_4 = 001_1111, "belongs to [m[+2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_01000 + 00_00000 + 01_00000 = 00_01000
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_0100 + 000_0000 + 000_0110 = 011_1010
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_0100 + 000_0000 + 111_1010 = 010_1110
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_01000 + 00_00000 + 11_00000 = 10_01000


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (00_01000 + 01_01111)_reduced_2_4 = 
(01_10111)_reduced_2_4 = 01_1011 >= 0, don't care.
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (011_1010 + 101_0111)_reduced_3_3 = 
(001_0001)_reduced_3_3 = 001_000 >= 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (010_1110 + 101_0111)_reduced_3_3 = 
(11_10111)_reduced_3_3 = 11_1011 < 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_01000 + 01_01111)_reduced_2_4 = 
(11_00000)_reduced_2_4 = 11_0000 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0101
q_neg = 0000

w[2] = 4 * w[1] - q[2] * D = 
1_11111010000111001110010001100000000 + 
0_00111111110101111111111100000000000 = 
0_00111001111101001110001101100000000

w[2] >= 0;
w[2]_reduced >> CLZ_D = 
00111001111101001110001101100000 >> 1 = 
00011100111110100111000110110000

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 11111101000011100111001000110000 = 4245582384
D[WIDTH-1:0] = 00111000000001010000000000100000 = 939851808
Q[WIDTH-1:0] = X / D = 4 = 00000000000000000000000000000010
REM[WIDTH-1:0] = 4245582384 - 939851808 * 4 = 486175152 = 00011100111110100111000110110000

CLZ_X = 0
CLZ_D = 2
CLZ_DIFF = CLZ_D - CLZ_X = 2
r_shift_num = CLZ_DIFF[0] = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(4 / 2) = 2;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11111101000011100111001000110000
Divisor[WIDTH-1:0] 		= 11100000000101000000000010000000

+ D = 0_11100000000101000000000010000000000
+2D = 1_11000000001010000000000100000000000
- D = 1_00011111111010111111111110000000000
-2D = 0_00111111110101111111111100000000000

根据D的值, 可得选择常数:
m[-1] = -22
m[ 0] = - 8
m[+1] = + 8
m[+2] = +22

// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0] = 0_00111111010000111001110010001100000

(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

w[1] = 4 * w[0] - q[1] * D = 
0_11111101000011100111001000110000000 + 
1_00011111111010111111111110000000000 = 
0_00011100111110100111000110110000000
(4 * w[1])_trunc_3_4 = 000_0111, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0100
q_neg = 0000

w[2] = 4 * w[1] - q[2] * D = 
0_01110011111010011100011011000000000 + 
0_00000000000000000000000000000000000 = 
0_01110011111010011100011011000000000

w[2] >= 0;
w[2]_reduced >> CLZ_D = 
01110011111010011100011011000000 >> 2 = 
00011100111110100111000110110000

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------





------------------------------------------------------------------------------------
ERROR FOUND:
dividend = 079aad02, divisor = 0000067f
opcode = 0
exp_quotient = 00012bab, exp_remainder = 0000012d, act_quotient = 00012baa, act_remainder = 000007ac
exp_divisor_is_zero = 0, dut_divisor_is_zero = 0
finished_test_num =   47847232, error_test_num =          1

------------------------------------------------------------------------------------
ERROR FOUND:
dividend = 3b92b337, divisor = 0000067f
opcode = 0
exp_quotient = 00092bac, exp_remainder = 000000e3, act_quotient = 00092ba9, act_remainder = 00000460
exp_divisor_is_zero = 0, dut_divisor_is_zero = 0

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00111011100100101011001100110111 = 999469879
D[WIDTH-1:0] = 00000000000000000000011001111111 = 1663
Q[WIDTH-1:0] = X / D = 601004 = 00000000000010010010101110101100
R[WIDTH-1:0] = 227 = 00000000000000000000000011100011

CLZ_X = 2
CLZ_D = 21
CLZ_DIFF = CLZ_D - CLZ_X = 19
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (20 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(21 / 2) = 11;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11101110010010101100110011011100
Divisor[WIDTH-1:0] 		= 11001111111000000000000000000000

+ D = 0_11001111111000000000000000000000000
+2D = 1_10011111110000000000000000000000000
- D = 1_00110000001000000000000000000000000
-2D = 0_01100000010000000000000000000000000
~ D = 1_00110000000111111111111111111111111
~2D = 0_01100000001111111111111111111111111

根据D的值, 可得选择常数:
m[-1] = -19
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

-m[-1]_reduced_2_5 = 01_00110
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 10_11100
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] = 0_00011101110010010101100110011011100
w_carry[0] = 0_00000000000000000000000000000000000
w[0] = 0_00011101110010010101100110011011100
(4 * w[0])_trunc_3_4 = 000_0111, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
w[1] = 4 * w[0] - q[1] * D = 
0_01110111001001010110011001101110000 + 
1_00110000001000000000000000000000000 = 
1_10100111010001010110011001101110000
(4 * w[1])_trunc_3_4 = 110_1001, "belongs to [-Inf, m[-1])" -> q[2] = -2
q_pos = 0100
q_neg = 0010

ITER[1]:
w[2] = 4 * w[1] - q[2] * D = 
0_10011101000101011001100110111000000 + 
1_10011111110000000000000000000000000 = 
0_00111100110101011001100110111000000
(4 * w[2])_trunc_3_4 = 000_1111, "belongs to [m[-1], m[0])" -> q[3] = +1
q_pos = 0100_01
q_neg = 0010_00

ITER[2]:
w[3] = 4 * w[2] - q[3] * D = 
0_11110011010101100110011011100000000 + 
1_00110000001000000000000000000000000 = 
0_00100011011101100110011011100000000
(4 * w[3])_trunc_3_4 = 000_1000, "belongs to [m[-1], m[0])" -> q[4] = +1
q_pos = 0100_0101
q_neg = 0010_0000

ITER[3]:
w[4] = 4 * w[3] - q[4] * D = 
0_10001101110110011001101110000000000 + 
1_00110000001000000000000000000000000 = 
1_10111101111110011001101110000000000
(4 * w[4])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[5] = -1
q_pos = 0100_0101_00
q_neg = 0010_0000_01

ITER[4]:
w[5] = 4 * w[4] - q[5] * D = 
0_11110111111001100110111000000000000 + 
0_11001111111000000000000000000000000 = 
1_11000111110001100110111000000000000
(4 * w[5])_trunc_3_4 = 111_0001, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0100_0101_0000
q_neg = 0010_0000_0101

ITER[5]:
w[6] = 4 * w[5] - q[6] * D = 
1_00011111000110011011100000000000000 + 
0_11001111111000000000000000000000000 = 
1_11101110111110011011100000000000000
(4 * w[5])_trunc_3_4 = 111_1011, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0100_0101_0000_00
q_neg = 0010_0000_0101_00



w_sum = 1c7c80ff8 = 0_00111000111110010000000111111111000
w_cry = c766b6008 = 1_10001110110011010110110000000001000
1_11000111110001100110111000000000000

temp[0] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 01_00110 = 01_10100
temp[1] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 000_0110 = 100_1100
temp[2] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 111_1010 = 100_0000
temp[3] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 10_11100 = 11_01010

+ D = 0_11001111111000000000000000000000000 -> 11_00111, 011_0011
(temp[0] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (01_10100 + 11_00111)_reduced_2_4 = 
(00_11011)_reduced_2_4 = 00_1101 >= 0
(temp[1] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_1100 + 011_0011)_reduced_3_3 = 
(111-1111)_reduced_3_3 = 111_111 < 0
(temp[2] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_0000 + 011_0011)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[3] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (11_01010 + 11_00111)_reduced_2_4 = 
(10_10001)_reduced_2_4 = 10_1000 < 0
根据比较结果(Sign Detection, SD)可得 -> q = -1 -> 又出错了









ITER[6]:
w[7] = 4 * w[6] - q[7] * D = 
1_10111011111001101110000000000000000 + 
0_00000000000000000000000000000000000 = 
1_10111011111001101110000000000000000
(4 * w[5])_trunc_3_4 = 110_1110, "belongs to [m[-1], m[0])" -> q[8] = -1
q_pos = 0100_0101_0000_0000
q_neg = 0010_0000_0101_0001


// ---------------------------------------------------------------------------------------------------------------------------------------





// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00011110011010101011100001011011 = 510310491
D[WIDTH-1:0] = 00000000000000000000011001111111 = 1663
Q[WIDTH-1:0] = X / D = 306861 = 00000000000001001010111010101101
R[WIDTH-1:0] = 648 = 00000000000000000000001010001000

CLZ_X = 3
CLZ_D = 21
CLZ_DIFF = CLZ_D - CLZ_X = 18
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (19 % 2) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(20 / 2) = 10;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11110011010101011100001011011000
Divisor[WIDTH-1:0] 		= 11001111111000000000000000000000

+ D = 0_11001111111000000000000000000000000
+2D = 1_10011111110000000000000000000000000
- D = 1_00110000001000000000000000000000000
-2D = 0_01100000010000000000000000000000000
~ D = 1_00110000000111111111111111111111111
~2D = 0_01100000001111111111111111111111111

根据D的值, 可得选择常数:
m[-1] = -19
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

-m[-1]_reduced_2_5 = 01_00110
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 10_11100
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] = 0_00111100110101010111000010110110000
w_carry[0] = 0_00000000000000000000000000000000000
w[0] = 0_00111100110101010111000010110110000
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
w[1] = 4 * w[0] - q[1] * D = 
0_11110011010101011100001011011000000 + 
1_00110000001000000000000000000000000 = 
0_00100011011101011100001011011000000
(4 * w[1])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0101
q_neg = 0000

ITER[1]:
w[2] = 4 * w[1] - q[2] * D = 
0_10001101110101110000101101100000000 + 
1_00110000001000000000000000000000000 = 
1_10111101111101110000101101100000000
(4 * w[2])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0101_00
q_neg = 0000_01

ITER[2]:
w[3] = 4 * w[2] - q[3] * D = 
0_11110111110111000010110110000000000 + 
0_11001111111000000000000000000000000 = 
1_11000111101111000010110110000000000
(4 * w[3])_trunc_3_4 = 111_0001, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0101_0000
q_neg = 0000_0101

ITER[3]:
w[4] = 4 * w[3] - q[4] * D = 
1_00011110111100001011011000000000000 + 
0_11001111111000000000000000000000000 = 
1_11101110110100001011011000000000000
(4 * w[4])_trunc_3_4 = 111_1011, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0101_0000_00
q_neg = 0000_0101_00


w_sum = 1c79e03f8 = 0_0011-10001-11100111100000001111111000
w_cry = c76436808 = 1_10001110110010000110110100000001000
1_11000111101111000010110110000000000 -> 00_01111, 100_0111

temp[0] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 01_00110 = 01_10100
temp[1] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 000_0110 = 100_1100
temp[2] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 111_1010 = 100_0000
temp[3] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 10_11100 = 11_01010

+ D = 0_11001111111000000000000000000000000 -> 11_00111, 011_0011
(temp[0] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (01_10100 + 11_00111)_reduced_2_4 = 
(00_11011)_reduced_2_4 = 00_1101 >= 0
(temp[1] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_1100 + 011_0011)_reduced_3_3 = 
(111_1111)_reduced_3_3 = 111_111 < 0
(temp[2] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_0000 + 011_0011)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[3] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (11_01010 + 11_00111)_reduced_2_4 = 
(10_10001)_reduced_2_4 = 10_1000 < 0
根据比较结果(Sign Detection, SD)可得 -> q = -1 -> 又出错了






// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000111100110101010110100000010 = 127577346
D[WIDTH-1:0] = 00000000000000000000011001111111 = 1663
Q[WIDTH-1:0] = X / D = 76715 = 00000000000000010010101110101011
R[WIDTH-1:0] = 301 = 00000000000000000000000100101101

CLZ_X = 5
CLZ_D = 21
CLZ_DIFF = CLZ_D - CLZ_X = 16
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (17 % 2) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(18 / 2) = 9;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11110011010101011010000001000000
Divisor[WIDTH-1:0] 		= 11001111111000000000000000000000

+ D = 0_11001111111000000000000000000000000
+2D = 1_10011111110000000000000000000000000
- D = 1_00110000001000000000000000000000000
-2D = 0_01100000010000000000000000000000000
~ D = 1_00110000000111111111111111111111111
~2D = 0_01100000001111111111111111111111111

根据D的值, 可得选择常数:
m[-1] = -19
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

-m[-1]_reduced_2_5 = 01_00110
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 10_11100

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// TODO
// 最后一次迭代的余数
w[final] = w[11];
w[11] = 4 * w[10] - q[11] * D = 
1_10010001010110000000000000000000000 + 
0_00000000000000000000000000000000000 = 
1_10010001010110000000000000000000000 < 0
// 最后一次迭代的商
q_pos = 0001_0101_0000_0100_0000_00
q_neg = 0000_0000_0110_0001_0101_00
corr(q_pos - q_neg) = 01010010100010101011

(10010001010110000000000000000000 + 11100000000100000000000000000000) >> 19 = 
01110001011010000000000000000000 >> 19 = 
00000000000000000000111000101101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] = 0_00111100110101010110100000010000000
w_carry[0] = 0_00000000000000000000000000000000000
w[0] = 0_00111100110101010110100000010000000
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
w[1] = 4 * w[0] - q[1] * D = 
0_11110011010101011010000001000000000 + 
1_00110000001000000000000000000000000 = 
0_00100011011101011010000001000000000
(4 * w[1])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0101
q_neg = 0000

ITER[1]:
w[2] = 4 * w[1] - q[2] * D = 
0_10001101110101101000000100000000000 + 
1_00110000001000000000000000000000000 = 
1_10111101111101101000000100000000000
(4 * w[2])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0101_00
q_neg = 0000_01

ITER[2]:
w[3] = 4 * w[2] - q[3] * D = 
0_11110111110110100000010000000000000 + 
0_11001111111000000000000000000000000 = 
1_11000111101110100000010000000000000
(4 * w[3])_trunc_3_4 = 111_0001, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0101_0000
q_neg = 0000_0101

ITER[3]:
w[4] = 4 * w[3] - q[4] * D = 
1_00011110111010000001000000000000000 + 
0_11001111111000000000000000000000000 = 
1_11101110110010000001000000000000000
(4 * w[4])_trunc_3_4 = 111_1011, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0101_0000_00
q_neg = 0000_0101_00

w_sum = 0b93e7fc0 = 0_00010111001001111100111111111000000
w_carry = ebd020040 = 1_11010111101000000100000000001000000
(4 * w_sum)_reduced_3_4 + (4 * w_carry)_reduced_3_4 = 
000_0101 + 111_0101 = 111_1010, , "belongs to [m[0], m[+1])" -> q[5] = 0
-> 这也不会造成q[5] = -1.....

// ---------------------------------------------------------------------------------------------------------------------------------------

w_sum_pre = 1c72fdff8 = 0_0011-1000111001011111101111111111000
w_carry_pre = c76a04008 = 1_1000-1110110101000000100000000001000
1_11000111101110100000010000000000000 -> 100_0111


temp[0] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 01_00110 = 01_10100
temp[1] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 000_0110 = 100_1100
temp[2] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1000 + 000_1110 + 111_1010 = 100_0000
temp[3] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_10001 + 00_11101 + 10_11100 = 11_01010

+ D = 0_11001111111000000000000000000000000 -> 11_00111, 011_0011
(temp[0] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (01_10100 + 11_00111)_reduced_2_4 = 
(00_11011)_reduced_2_4 = 00_1101 >= 0
(temp[1] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_1100 + 011_0011)_reduced_3_3 = 
(111_1111)_reduced_3_3 = 111_111 < 0
(temp[2] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (100_0000 + 011_0011)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[3] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (11_01010 + 11_00111)_reduced_2_4 = 
(10_10001)_reduced_2_4 = 10_1000 < 0
根据比较结果(Sign Detection, SD)可得 -> q = -1 -> 又出错了


// ---------------------------------------------------------------------------------------------------------------------------------------










ITER[4]:
w[5] = 4 * w[4] - q[5] * D = 
1_10111011001000000100000000000000000 + 
0_00000000000000000000000000000000000 = 
1_10111011001000000100000000000000000
(4 * w[5])_trunc_3_4 = 110_1110, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0101_0000_0000
q_neg = 0000_0101_0001


ITER[5]:
w[6] = 4 * w[5] - q[6] * D = 
0_11101100100000010000000000000000000 + 
0_11001111111000000000000000000000000 = 
1_10111100011000010000000000000000000
(4 * w[6])_trunc_3_4 = 110_1111, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0101_0000_0000_00
q_neg = 0000_0101_0001_01

ITER[6]:
w[7] = 4 * w[6] - q[7] * D = 
0_11110001100001000000000000000000000 + 
0_11001111111000000000000000000000000 = 
1_11000001011001000000000000000000000
(4 * w[7])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[8] = -1
q_pos = 0101_0000_0000_0000
q_neg = 0000_0101_0001_0101

ITER[7]:
w[8] = 4 * w[7] - q[8] * D = 
1_00000101100100000000000000000000000 + 
0_11001111111000000000000000000000000 = 
1_11010101011100000000000000000000000
(4 * w[8])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[9] = -1
q_pos = 0101_0000_0000_0000_00
q_neg = 0000_0101_0001_0101_01

// TODO
ITER[8]:
w[9] = 4 * w[8] - q[9] * D = 
0_11111000111101100000000000000000000 + 
0_11001000000000000000000000000000000 = 
1_11000000111101100000000000000000000
(4 * w[9])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[10] = -1
q_pos = 0001_0101_0110_0000_0000
q_neg = 0000_0000_0000_1000_0101

ITER[9]:
w[10] = 4 * w[9] - q[10] * D = 
1_00000011110110000000000000000000000 + 
0_11001000000000000000000000000000000 = 
1_11001011110110000000000000000000000
(4 * w[10])_trunc_3_4 = 111_0010, "belongs to [m[-1], m[0])" -> q[11] = -1
q_pos = 0001_0101_0110_0000_0000_00
q_neg = 0000_0000_0000_1000_0101_01

ITER[10]:
w[11] = 4 * w[10] - q[11] * D = 
1_00101111011000000000000000000000000 + 
0_11001000000000000000000000000000000 = 
1_11110111011000000000000000000000000
(4 * w[11])_trunc_3_4 = 111_1101, "belongs to [m[0], m[+1])" -> q[12] = 0
q_pos = 0001_0101_0110_0000_0000_0000
q_neg = 0000_0000_0000_1000_0101_0100

ITER[11]:
w[12] = 4 * w[11] - q[12] * D = 
1_11011101100000000000000000000000000 + 
0_00000000000000000000000000000000000 = 
1_11011101100000000000000000000000000
(4 * w[12])_trunc_3_4 = 111_0111, "belongs to [m[-1], m[0])" -> q[13] = -1
q_pos = 0001_0101_0110_0000_0000_0000_00
q_neg = 0000_0000_0000_1000_0101_0100_01

ITER[12]:
w[13] = 4 * w[12] - q[13] * D = 
1_01110110000000000000000000000000000 + 
0_11001000000000000000000000000000000 = 
0_00111110000000000000000000000000000
(4 * w[13])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[14] = +1
q_pos = 0001_0101_0110_0000_0000_0000_0001
q_neg = 0000_0000_0000_1000_0101_0100_0100

w[14] = 4 * w[13] - q[14] * D = 
0_11111000000000000000000000000000000 + 
1_00111000000000000000000000000000000 = 
0_00110000000000000000000000000000000 >= 0


corr(q_pos - q_neg) = 0001010101010111101010111101





// ---------------------------------------------------------------------------------------------------------------------------------------









if(q[6] = +1) begin
ITER[4]:
w[5] = 4 * w[4] - q[5] * D = 
1_00010001111110001111011000000000000 + 
1_00111000000000000000000000000000000 = 
0_01001001111110001111011000000000000
(4 * w[5])_trunc_3_4 = 001_0010 -> q[6] = +1
q_pos = 0001_0101_0101
q_neg = 0000_0000_0000

ITER[5]:
w[6] = 4 * w[5] - q[6] * D = 
1_00100111111000111101100000000000000 + 
1_00111000000000000000000000000000000 = 
0_01011111111000111101100000000000000
(4 * w[6])_trunc_3_4 = 001_0111, "belongs to [m[+2], +Inf)" -> q[7] = +2
q_pos = 0001_0101_0101_10
q_neg = 0000_0000_0000_00

ITER[6]:
w[7] = 4 * w[6] - q[7] * D = 
1_01111111100011110110000000000000000 + 
0_01110000000000000000000000000000000 = 
1_11101111100011110110000000000000000
(4 * w[7])_trunc_3_4 = 111_1011, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0001_0101_0101_1000
q_neg = 0000_0000_0000_0000

w_sum_pre = f0f3ec007 = 1_11100001111001111101100000000000111
w_carry_pre = 3efdffff9 = 0_01111101111110111111111111111111001
0_01011111111000111101100000000000000
-2D = 0_01110000000000000000000000000000000 -> 01_11000, 001_1100
~2D = 0_01101111111111111111111111111111111 -> 01_10111, 001_1011
使用~2D
temp[0] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_00011 + 11_11011 + 01_00110 = 11_00100
temp[1] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_0001 + 111_1101 + 000_0110 = 110_0100
temp[2] = ((16 * w_sum)_reduced_3_4 + (16 * w_carry)_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_0001 + 111_1101 + 111_1010 = 101_1000
temp[3] = ((16 * w_sum)_reduced_2_5 + (16 * w_carry)_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_00011 + 11_11011 + 10_11100 = 00_11010


(temp[0] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (11_00100 + 01_10111)_reduced_2_4 = 
(00_11011)_reduced_2_4 = 00_1101 >= 0
(temp[1] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (110_0100 + 001_1011)_reduced_3_3 = 
(111_1111)_reduced_3_3 = 111_111 < 0
(temp[2] + (-4 * q * D)_reduced_3_4)_reduced_3_3 = (101_1000 + 001_1011)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[3] + (-4 * q * D)_reduced_2_5)_reduced_2_4 = (00_11010 + 01_10111)_reduced_2_4 = 
(10_10001)_reduced_2_4 = 10_1000 < 0, don't care.
根据比较结果(Sign Detection, SD)可得 -> q = -1 


if(q[8] = -1) begin
ITER[7]:
w[8] = 4 * w[7] - q[8] * D = 
1_10111110001111011000000000000000000 + 
0_11001000000000000000000000000000000 = 
0_10000110001111011000000000000000000 -> 溢出, 错误
end





















测试初始化操作

指数是奇数:
a_frac = 1.1010001111
a_frac << 1 = 11.0100011110
sqrt(a_frac << 1) = 1.11001111100101100000010110001101011001111111111011
a_frac >> 1 = 0.11010001111


r_s[0] = 1 - (a_frac >> 1) = 11_11010001111000
r_c[0] = 00_00000000000000
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

a_frac[9] = 1, s[1] = 0
-> 
r_s[1] = 11_01000111100000
r_c[1] = 00_00000000000000
rt_pos  = 01_00
rt_neg  = 00_00
rt[1]   = 01_00
rt_m[1] = 00_11

r[1] = r_s[1] + r_c[1] = 
11_01000111100000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_11
11_01000111100000 + 
01_11000000000000 = 
01_00000111100000


a_frac << 1 = 11.0100011110
sqrt(a_frac << 1) = 1.11001111100101100000010110001101011001111111111011
rt_real = 1.1
rt_real ^ 2 = 10.01000000000000000000000000000000000000000000000000
rem_real = 11.0100011110 - 10.01000000000000000000000000000000000000000000000000 = 
1.00000111100000000000000000000000000000000000000000
// r[1] is correct


// ================================================================================================================================================
指数是奇数:
a_frac = 1.0010111001
a_frac << 1 = 10.0101110010
sqrt(a_frac << 1) = 1.10001001011000101010001101111111110011110000111001
a_frac >> 1 = 0.10010111001

r_s[0] = 1 - (a_frac >> 1) = 11_10010111001000
r_c[0] = 00_00000000000000
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

a_frac[9] = 0, s[1] = -1
-> 
r_s[1] = 10_01011100100000
r_c[1] = 01_11000000000000
rt_pos  = 01_00
rt_neg  = 00_01
rt[1]   = 00_11
rt_m[1] = 00_10

r[1] = r_s[1] + r_c[1] = 
00_00011100100000

a_frac << 1 = 10.0101110010
sqrt(a_frac << 1) = 1.10001001011000101010001101111111110011110000111001
rt_real = 1.1
rt_real ^ 2 = 10.01000000000000000000000000000000000000000000000000
rem_real = 10.0101110010 - 10.01000000000000000000000000000000000000000000000000 = 
0.00011100100000000000000000000000000000000000000000
// r[1] is correct

// ================================================================================================================================================
指数是偶数:
a_frac = 1.1010111110
sqrt(a_frac) = 1.01001100010111000111101011010100100111101111000000
a_frac >> 2 = 0.011010111110

r_s[0] = 1 - (a_frac >> 2) = 11_01101011111000
r_c[0] = 00_00000000000000
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

a_frac[9] = 1, s[1] = -1
-> 
r_s[1] = 01_10101111100000
r_c[1] = 01_11000000000000
rt_pos  = 01_00
rt_neg  = 00_01
rt[1]   = 00_11
rt_m[1] = 00_10

r[1] = r_s[1] + r_c[1] = 
11_01101111100000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_11
11_01101111100000 + 
01_11000000000000 = 
01_00101111100000


a_frac = 1.1010111110
sqrt(a_frac) = 1.01001100010111000111101011010100100111101111000000
rt_real = 1.0
rt_real ^ 2 = 1.00000000000000000000000000000000000000000000000000
rem_real = 1.1010111110 - 1.00000000000000000000000000000000000000000000000000 = 
0.10101111100000000000000000000000000000000000000000
// r[1] is correct


// ================================================================================================================================================
指数是偶数:
a_frac = 1.0011100101
sqrt(a_frac) = 1.00011011001011101001001001010100100111100100011111
a_frac >> 2 = 0.010011100101

r_s[0] = 1 - (a_frac >> 2) = 11_01001110010100
r_c[0] = 00_00000000000000
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

a_frac[9] = 0, s[1] = -2
-> 
r_s[1] = 01_00111001010000
r_c[1] = 11_00000000000000
rt_pos  = 01_00
rt_neg  = 00_10
rt[1]   = 00_10
rt_m[1] = 00_01

r[1] = r_s[1] + r_c[1] = 
00_00111001010000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_11
11_01101111100000 + 
01_11000000000000 = 
01_00101111100000


a_frac = 1.0011100101
sqrt(a_frac) = 1.00011011001011101001001001010100100111100100011111
rt_real = 1.0
rt_real ^ 2 = 1.00000000000000000000000000000000000000000000000000
rem_real = 1.0011100101 - 1.00000000000000000000000000000000000000000000000000 = 
0.00111001010000000000000000000000000000000000000000
// r[1] is correct









// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00100010100001110000011111001110 = 579274702
D[WIDTH-1:0] = 00100101000011111110100011000110 = 621799622
Q[WIDTH-1:0] = X / D = 0 = 00000000000000000000000000000000
REM[WIDTH-1:0] = 579274702 - 621799622 * 0 = 579274702 = 00100010100001110000011111001110

CLZ_X = 0
CLZ_D = 0
CLZ_DIFF = CLZ_D - CLZ_X = 0
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (0 % 4) = 3;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(1 / 4) = 1;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 10001010000111000001111100111000
Divisor[WIDTH-1:0] 		= 10010100001111111010001100011000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_0010100001111111010001100011000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_0101000011111110100011000110000000
~ D[(WIDTH + 1 + log2(N))-1:0] = 110_1101011110000000101110011100111111
- D[(WIDTH + 1 + log2(N))-1:0] = 110_1101011110000000101110011101000000
~2D[(WIDTH + 1 + log2(N))-1:0] = 101_1010111100000001011100111001111111
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_1010111100000001011100111010000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[4] = 101_1000011001110011011001000010000000 < 0;
(w[final] / 2) + (D) = 110_1100001100111001101100100001000000 + 001_0010100001111111010001100011000000 = 
111_1110101110111000111110000100000000 < 0 -> (w[final] / 2) "belongs to [-2D, -D)";
// 最后一次迭代的商
q_pos = 1000
q_neg = 0110

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 0010;
(w[final] / 2) "belongs to [-2D, -D)" -> quotient_correction_coefficient = -2;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 0000;

(w[final] / 2) "belongs to [-2D, -D)" -> remainder_correction_coefficient = -2;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
(110_1100001100111001101100100001000000 + 010_0101000011111110100011000110000000) >> 2 = 
10001010000111000001111100111000 >> 2 = 
00100010100001110000011111001110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_0010001010000111000001111100111000
w_sum_translation[0] = w_sum[0] =  000_0010001010000111000001111100111000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_0000000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_1110101000001111011111000000001110
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_0000101000000000000001110011100010
w_sum_translation[1] = 111_1110101000001111011111000000001110
w_carry_translation[1] = 110_0000101000000000000001110011100010
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_10 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_0010001010000111000001111100111000 +
	110_1101011110000000101110011101000000
) = 2 * 110_1111101000000111110000011001111000 = 
101_1111010000001111100000110011110000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_1001000011100000011110100001011000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_1010100000111101000110001100001000
w_sum_translation[2] = 111_1001000011100000011110100001011000
w_carry_translation[2] = 110_1010100000111101000110001100001000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 11_10 -> q[3] = -1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	101_1111010000001111100000110011110000 +
	001_0010100001111111010001100011000000
) = 2 * 111_0001110010001110110010010110110000 = 
110_0011100100011101100100101101100000
q_pos = 100
q_neg = 011

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_0010000101000100010010011100100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_1010000111110101011010000100100000
w_sum_translation[3] = 000_0010000101000100010010011100100000
w_carry_translation[3] = 110_1010000111110101011010000100100000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	110_0011100100011101100100101101100000 +
	001_0010100001111111010001100011000000
) = 2 * 111_0110000110011100110110010000100000 = 
110_1100001100111001101100100001000000
q_pos = 1000
q_neg = 0110

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_0100001010001000100100111001000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
101_0100001111101010110100001001000000
w_sum_translation[4] = 110_0100001010001000100100111001000000
w_carry_translation[4] = 111_0100001111101010110100001001000000
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	110_1100001100111001101100100001000000 +
	000_0000000000000000000000000000000000
) = 2 * 110_1100001100111001101100100001000000 = 
101_1000011001110011011001000010000000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00111011010100000000101001100101 = 995101285
D[WIDTH-1:0] = 00110001000001110111101100111010 = 822573882
Q[WIDTH-1:0] = X / D = 1 = 00000000000000000000000000000001
REM[WIDTH-1:0] = 995101285 - 822573882 * 1 = 172527403 = 00001010010010001000111100101011

CLZ_X = 2
CLZ_D = 2
CLZ_DIFF = CLZ_D - CLZ_X = 0
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (0 % 4) = 3;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(1 / 4) = 1;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 11101101010000000010100110010100
Divisor[WIDTH-1:0] 		= 11000100000111011110110011101000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_1000100000111011110110011101000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 011_0001000001110111101100111010000000
~ D[(WIDTH + 1 + log2(N))-1:0] = 110_0111011111000100001001100010111111
- D[(WIDTH + 1 + log2(N))-1:0] = 110_0111011111000100001001100011000000
~2D[(WIDTH + 1 + log2(N))-1:0] = 100_1110111110001000010011000101111111
-2D[(WIDTH + 1 + log2(N))-1:0] = 100_1110111110001000010011000110000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[4] = 000_1010010010001000111100101011000000 >= 0;
(w[final] / 2) + (-D) = 000_0101001001000100011110010101100000 + 110_0111011111000100001001100011000000 = 
110_1100101000001000100111111000100000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1010
q_neg = 1001

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 0001;
(w[final] / 2) "belongs to [-2D, -D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 0001;

(w[final] / 2) "belongs to [-2D, -D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
00101001001000100011110010101100 >> 2 = 
00001010010010001000111100101011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_0011101101010000000010100110010100
w_sum_translation[0] = w_sum[0] =  000_0011101101010000000010100110010100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_0000000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_1001100100101000010110001001010110
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_1100110100000000000010001001010010
w_sum_translation[1] = 110_1001100100101000010110001001010110
w_carry_translation[1] = 110_1100110100000000000010001001010010
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_10 -> q[2] = -2
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_0011101101010000000010100110010100 +
	110_0111011111000100001001100011000000
) = 2 * 110_1011001100010100001100001001010100 = 
101_0110011000101000011000010010101000
q_pos = 10
q_neg = 10

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
010_1000100010111111110001110100001000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_0110010010000000011000100101001000
w_sum_translation[2] = 000_1000100010111111110001110100001000
w_carry_translation[2] = 000_0110010010000000011000100101001000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_00 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	101_0110011000101000011000010010101000 +
	011_0001000001110111101100111010000000
) = 2 * 000_0111011010100000000101001100101000 = 
000_1110110101000000001010011001010000
q_pos = 101
q_neg = 100

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
101_0011011111110111000001100111111110
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
001_1001001000010001100110010000100010
w_sum_translation[3] = 111_0011011111110111000001100111111110
w_carry_translation[3] = 111_1001001000010001100110010000100010
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_11 -> q[4] = -1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_1110110101000000001010011001010000 +
	110_0111011111000100001001100011000000
) = 2 * 111_0110010100000100010011111100010000 = 
110_1100101000001000100111111000100000
q_pos = 1010
q_neg = 1001

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
010_0101101110111010100011010100111000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_0100100011001110011001010110001000
w_sum_translation[4] = 000_0101101110111010100011010100111000
w_carry_translation[4] = 000_0100100011001110011001010110001000
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	110_1100101000001000100111111000100000 +
	001_1000100000111011110110011101000000
) = 2 * 000_0101001001000100011110010101100000 = 
000_1010010010001000111100101011000000



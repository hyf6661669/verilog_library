尝试的记录，无效.

接"test_1.sv"
选择函数来自于参考论文的"Fig. 6 (c)":
case(w_sum[i][MSB-1:MSB-2], w_carry[i][MSB-1:MSB-2])
	4'b00_00:	q[i+1] = +1;
	4'b00_01:	q[i+1] = +1;
	4'b00_10:	q[i+1] = +0;
	4'b00_11:	q[i+1] = +0;
	4'b01_00:	q[i+1] = +1;
	4'b01_01:	q[i+1] = +2;
	4'b01_10:	q[i+1] = +0;
	4'b01_11:	q[i+1] = +0;
	4'b10_00:	q[i+1] = -0;
	4'b10_01:	q[i+1] = -0;
	4'b10_10:	q[i+1] = -2;
	4'b10_11:	q[i+1] = -1;
	4'b11_00:	q[i+1] = -0;
	4'b11_01:	q[i+1] = -0;
	4'b11_10:	q[i+1] = -1;
	4'b11_11:	q[i+1] = -1;
endcase

// 注意: 后面发现这个改变没卵用...
对于最后一次迭代，尝试使用新的特别选择函数, 其实不是最后一次迭代也能使用下面这个选择函数.
case(w_sum[i][MSB-1:MSB-2], w_carry[i][MSB-1:MSB-2], q[i])
	4'b00_00:	q[i+1] = +1;
	4'b00_01:	q[i+1] = (q[i] > 0) ? +2: +1;
	4'b00_10:	q[i+1] = +0;
	4'b00_11:	q[i+1] = +0;
	4'b01_00:	q[i+1] = (q[i] > 0) ? +2: +1;
	4'b01_01:	q[i+1] = +2;
	4'b01_10:	q[i+1] = +0;
	4'b01_11:	q[i+1] = +0;
	4'b10_00:	q[i+1] = -0;
	4'b10_01:	q[i+1] = -0;
	4'b10_10:	q[i+1] = -2;
	4'b10_11:	q[i+1] = (q[i] < 0) ? -2: -1;
	4'b11_00:	q[i+1] = -0;
	4'b11_01:	q[i+1] = -0;
	4'b11_10:	q[i+1] = (q[i] < 0) ? -2: -1;
	4'b11_11:	q[i+1] = -1;
endcase


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000010000000110000 = 8240
Q[WIDTH-1:0] = X / D = 87 = 000000000000000001010111
REM[WIDTH-1:0] = 717047 - 8240 * 87 = 167 = 000000000000000010100111

CLZ_X = 4
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 6
迭代次数
iter_num = CLZ_DIFF + 1 + 1 = 8
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101011110000111101110000
Divisor[WIDTH-1:0] 		= 100000001100000000000000

+ D[(WIDTH + 2)-1:0] = 001_00000001100000000000000
+2D[(WIDTH + 2)-1:0] = 010_00000011000000000000000
- D[(WIDTH + 2)-1:0] = 110_11111110100000000000000
-2D[(WIDTH + 2)-1:0] = 101_11111101000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次按照特殊的选择函数来选
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +2
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	011_00001001101110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000110101110000000000 = 
010_00001101011100000000000
q_pos = 1010_1110
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
100_00100000111000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
011_11110100000000000000000
w_sum_translation[8] = 110_00100000111000000000000
w_carry_translation[8] = 001_11110100000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_01 -> q[9] = 0
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_00001101011100000000000 +
	101_11111101000000000000000
) = 2 * 000_00001010011100000000000 = 
000_00010100111000000000000
// 最后一次迭代的余数
w[final] = w[8];
w[final] = 000_00010100111000000000000 >= 0
// 最后一次迭代的商
q[8] = +1
q_pos = 1010_1110
q_neg = 0000_0000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
10101110
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 1010111
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
000000101001110000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
000000101001110000000000 >> 10 = 
000000000000000010100111

// 不改变QDS
q[7] = +2
q[8] = +1
q_pos = 1010_1101
q_neg = 0000_0000
w[final] = w[8];
w[final] = 010_00010111111000000000000 >= 0

q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
10101101
q_calculated = (q_calculated_pre[(WIDTH + 1) - 1:0] + 1) >> 1 = 1010111
w[final] / 2 =  = 001_00001011111100000000000
001_00001011111100000000000 + (-D) = 
001_00001011111100000000000 + 110_11111110100000000000000 = 000_00001010011100000000000
000_00001010011100000000000 >> (CLZ_D + 1) = 
000001010011100000000000 >> 11 = 
000000000000000010100111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000001000000011 = 515
Q[WIDTH-1:0] = X / D = 1392 = 000000000000010101110000
REM[WIDTH-1:0] = 717047 - 515 * 1392 = 167 = 000000000000000010100111

CLZ_X = 4
CLZ_D = 14
CLZ_DIFF = CLZ_D - CLZ_X = 10
迭代次数
iter_num = CLZ_DIFF + 1 + 1 = 12
// 最后一次按照特殊的选择函数来选
w_sum_translation[11] = 000_11110000000000000000000
w_carry_translation[11] = 001_10111010000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 00_01 -> q[12] = +2
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	010_01010110100000000000000 +
	110_11111110100000000000000
) = 2 * 001_01010101000000000000000 = 
010_10101010000000000000000
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	010_10101010000000000000000 +
	101_11111101000000000000000
) = 2 * 000_10100111000000000000000 = 
001_01001110000000000000000
// 最后一次迭代的余数
w[final] = w[12];
w[final] = 001_01001110000000000000000 >= 0
// 最后一次迭代的商
q[12] = +1
q_pos = 1010_1110_0000
q_neg = 0000_0000_0000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
101011100000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 10101110000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
001010011100000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
001010011100000000000000 >> 14 = 
000000000000000010100111

// 不改变QDS
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	010_01010110100000000000000 +
	110_11111110100000000000000
) = 2 * 001_01010101000000000000000 = 
010_10101010000000000000000
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	010_10101010000000000000000 +
	110_11111110100000000000000
) = 2 * 001_10101000100000000000000 = 
011_01010001000000000000000

w[final] = w[12] = 011_01010001000000000000000 >= 0
q[11] = +1
q[12] = +1
q_pos = 1010_1101_1111
q_neg = 0000_0000_0000
q_pos - q_neg = 101011011111
q_calculated = (101011011111 + 1) >> 1 = 10101110000

011_01010001000000000000000 / 2 = 001_10101000100000000000000
001_10101000100000000000000 + (-D) = 
001_10101000100000000000000 + 110_11111110100000000000000 = 000_10100111000000000000000
000_10100111000000000000000 >> (CLZ_D + 1) = 
010100111000000000000000 >> 15 = 
000000000000000010100111

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 2)-1:0] =  001_01011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_10111100001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11111101000000000000000
w_sum_translation[1] = 000_10111100001111011100000
w_carry_translation[1] = 111_11111101000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01011110000111101110000 +
	110_11111110100000000000000
) = 2 * 000_01011100100111101110000 = 
000_10111001001111011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_01111000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11111010000000000000000
w_sum_translation[2] = 001_01111000011110111000000
w_carry_translation[2] = 111_11111010000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_10111001001111011100000 +
	000_00000000000000000000000
) = 2 * 000_10111001001111011100000 = 
001_01110010011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_11110000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_11110100000000000000000
w_sum_translation[3] = 000_11110000111101110000000
w_carry_translation[3] = 001_11110100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_01 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_01110010011110111000000 +
	000_00000000000000000000000
) = 2 * 001_01110010011110111000000 = 
010_11100100111101110000000
q_pos = 1001
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_11110100111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11010010000000000000000
w_sum_translation[4] = 001_11110100111011100000000
w_carry_translation[4] = 001_11010010000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[5] = +2
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	010_11100100111101110000000 +
	110_11111110100000000000000
) = 2 * 001_11100011011101110000000 = 
011_11000110111011100000000
q_pos = 1010_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_10110111110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11010000000000000000000
w_sum_translation[5] = 001_10110111110111000000000
w_carry_translation[5] = 001_11010000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	011_11000110111011100000000 +
	101_11111101000000000000000
) = 2 * 001_11000011111011100000000 = 
011_10000111110111000000000
q_pos = 1010_10
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_00110101101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_11010100000000000000000
w_sum_translation[6] = 001_00110101101110000000000
w_carry_translation[6] = 001_11010100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_01 -> q[7] = +2
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_10000111110111000000000 +
	101_11111101000000000000000
) = 2 * 001_10000100110111000000000 = 
011_00001001101110000000000
q_pos = 1010_110
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_00111001011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_11010100000000000000000
w_sum_translation[7] = 000_00111001011100000000000
w_carry_translation[7] = 001_11010100000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	011_00001001101110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000110101110000000000 = 
010_00001101011100000000000
q_pos = 1010_1101
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
110_00100111111000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
011_11110000000000000000000
w_sum_translation[8] = 000_00100111111000000000000
w_carry_translation[8] = 001_11110000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 00_01 -> q[9] = +1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_00001101011100000000000 +
	110_11111110100000000000000
) = 2 * 001_00001011111100000000000 = 
010_00010111111000000000000
q_pos = 1010_1101_1
q_neg = 0000_0000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_01010010110000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
011_11011010000000000000000
w_sum_translation[9] = 000_01010010110000000000000
w_carry_translation[9] = 001_11011010000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_01 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	010_00010111111000000000000 +
	110_11111110100000000000000
) = 2 * 001_00010110011000000000000 = 
010_00101100110000000000000
q_pos = 1010_1101_11
q_neg = 0000_0000_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
110_11101100100000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
011_01101010000000000000000
w_sum_translation[10] = 000_11101100100000000000000
w_carry_translation[10] = 001_01101010000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 00_01 -> q[11] = +1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	010_00101100110000000000000 +
	110_11111110100000000000000
) = 2 * 001_00101011010000000000000 = 
010_01010110100000000000000
q_pos = 1010_1101_111
q_neg = 0000_0000_000

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
110_11110000000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
011_10111010000000000000000
w_sum_translation[11] = 000_11110000000000000000000
w_carry_translation[11] = 001_10111010000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 00_01 -> q[12] = +1
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	010_01010110100000000000000 +
	110_11111110100000000000000
) = 2 * 001_01010101000000000000000 = 
010_10101010000000000000000
q_pos = 1010_1101_1111
q_neg = 0000_0000_0000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000111011110000111101110 = 1958382
D[WIDTH-1:0] = 000000000000001110110100 = 948
Q[WIDTH-1:0] = X / D = 2065 = 000000000000100000010001
REM[WIDTH-1:0] = 1958382 - 948 * 2065 = 762 = 000000000000001011111010

CLZ_X = 3
CLZ_D = 14
CLZ_DIFF = CLZ_D - CLZ_X = 11
迭代次数
iter_num = CLZ_DIFF + 1 + 1 = 13
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111011110000111101110000
Divisor[WIDTH-1:0] 		= 111011010000000000000000

+ D[(WIDTH + 2)-1:0] = 001_11011010000000000000000
+2D[(WIDTH + 2)-1:0] = 011_10110100000000000000000
- D[(WIDTH + 2)-1:0] = 110_00100110000000000000000
-2D[(WIDTH + 2)-1:0] = 100_01001100000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[13];
w[final] = 110_10001100000000000000000 < 0
// 最后一次迭代的商
q[13] = 0
q_pos = 1000_0010_0100_0
q_neg = 0000_0001_0010_0
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
0001000000100100
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 000100000010001
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
110100011000000000000000 + 111011010000000000000000 = 
101111101000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
101111101000000000000000 >> 14 = 
000000000000001011111010
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000111011110000111101110 = 1958382
D[WIDTH-1:0] = 000000000111011010000000 = 30336
Q[WIDTH-1:0] = X / D = 64 = 0000000000000000000001000000
REM[WIDTH-1:0] = 1958382 - 30336 * 64 = 16878 = 0000000000000100000111101110

CLZ_X = 3
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 6
迭代次数
iter_num = CLZ_DIFF + 1 + 1 = 8
// 最后一次迭代的余数
w[final] = w[8];
w[final] = 100_10110110111000000000000 < 0
// 最后一次迭代的商
q[8] = +2
q_pos = 1000_0010
q_neg = 0000_0000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
10000010
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 1000000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
100101101101110000000000 + 111011010000000000000000 = 
100000111101110000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
100000111101110000000000 >> 9 = 
000000000100000111101110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_11011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_11011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_10111100001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_01001100000000000000000
w_sum_translation[1] = 001_10111100001111011100000
w_carry_translation[1] = 110_01001100000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11011110000111101110000 +
	110_00100110000000000000000
) = 2 * 000_00000100000111101110000 = 
000_00001000001111011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_01111000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_10011000000000000000000
w_sum_translation[2] = 001_01111000011110111000000
w_carry_translation[2] = 110_10011000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_00001000001111011100000 +
	000_00000000000000000000000
) = 2 * 000_00001000001111011100000 = 
000_00010000011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_11110000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
101_00110000000000000000000
w_sum_translation[3] = 000_11110000111101110000000
w_carry_translation[3] = 111_00110000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00010000011110111000000 +
	000_00000000000000000000000
) = 2 * 000_00010000011110111000000 = 
000_00100000111101110000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_11100001111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_01100000000000000000000
w_sum_translation[4] = 001_11100001111011100000000
w_carry_translation[4] = 110_01100000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00100000111101110000000 +
	000_00000000000000000000000
) = 2 * 000_00100000111101110000000 = 
000_01000001111011100000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11000011110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_11000000000000000000000
w_sum_translation[5] = 001_11000011110111000000000
w_carry_translation[5] = 110_11000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_01000001111011100000000 +
	000_00000000000000000000000
) = 2 * 000_01000001111011100000000 = 
000_10000011110111000000000
q_pos = 1000_00
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_10000111101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_10000000000000000000000
w_sum_translation[6] = 001_10000111101110000000000
w_carry_translation[6] = 111_10000000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_11 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_10000011110111000000000 +
	000_00000000000000000000000
) = 2 * 000_10000011110111000000000 = 
001_00000111101110000000000
q_pos = 1000_000
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_00001111011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_00000000000000000000000
w_sum_translation[7] = 001_00001111011100000000000
w_carry_translation[7] = 001_00000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 01_01 -> q[8] = +2
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	001_00000111101110000000000 +
	000_00000000000000000000000
) = 2 * 001_00000111101110000000000 = 
010_00001111011100000000000
q_pos = 1000_0010
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
100_10000110111000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
000_00110000000000000000000
w_sum_translation[8] = 110_10000110111000000000000
w_carry_translation[8] = 110_00110000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_10 -> q[9] = -2
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_00001111011100000000000 +
	100_01001100000000000000000
) = 2 * 110_01011011011100000000000 = 
100_10110110111000000000000
q_pos = 1000_0010_0
q_neg = 0000_0001_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
010_00000101110000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_11010000000000000000000
w_sum_translation[9] = 000_00000101110000000000000
w_carry_translation[9] = 000_11010000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_00 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	100_10110110111000000000000 +
	011_10110100000000000000000
) = 2 * 000_01101010111000000000000 = 
000_11010101110000000000000
q_pos = 1000_0010_01
q_neg = 0000_0001_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
101_11100111100000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
000_00010000000000000000000
w_sum_translation[10] = 111_11100111100000000000000
w_carry_translation[10] = 110_00010000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 11_10 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	000_11010101110000000000000 +
	110_00100110000000000000000
) = 2 * 110_11111011110000000000000 = 
101_11110111100000000000000
q_pos = 1000_0010_010
q_neg = 0000_0001_001

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
000_01011011000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
111_01001000000000000000000
w_sum_translation[11] = 000_01011011000000000000000
w_carry_translation[11] = 111_01001000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 00_11 -> q[12] = 0
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	101_11110111100000000000000 +
	001_11011010000000000000000
) = 2 * 111_11010001100000000000000 = 
111_10100011000000000000000
q_pos = 1000_0010_0100
q_neg = 0000_0001_0010

w_sum[12] = 2 * csa_sum(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
000_10110110000000000000000
w_carry[12] = 2 * csa_carry(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
110_10010000000000000000000
w_sum_translation[12] = 000_10110110000000000000000
w_carry_translation[12] = 110_10010000000000000000000
{w_sum_translation[12][MSB-1:MSB-2], w_carry_translation[12][MSB-1:MSB-2]} = 00_10 -> q[13] = 0
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	111_10100011000000000000000 +
	000_00000000000000000000000
) = 2 * 111_10100011000000000000000 = 
111_01000110000000000000000
q_pos = 1000_0010_0100_0
q_neg = 0000_0001_0010_0

w_sum[13] = 2 * csa_sum(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
001_01101100000000000000000
w_carry[13] = 2 * csa_carry(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
101_00100000000000000000000
w_sum_translation[13] = 111_01101100000000000000000
w_carry_translation[13] = 111_00100000000000000000000
{w_sum_translation[13][MSB-1:MSB-2], w_carry_translation[13][MSB-1:MSB-2]} = 11_11 -> q[14] = -1
w[13] = 2 * (w[12] - q[13] * D) = 2 * (
	111_01000110000000000000000 +
	000_00000000000000000000000
) = 2 * 111_01000110000000000000000 = 
110_10001100000000000000000
q_pos = 1000_0010_0100_00
q_neg = 0000_0001_0010_01

w_sum[14] = 2 * csa_sum(w_sum_translation[13], w_carry_translation[13], -q[14] * D) = 
011_00101100000000000000000
w_carry[14] = 2 * csa_carry(w_sum_translation[13], w_carry_translation[13], -q[14] * D) = 
101_10100000000000000000000
w_sum_translation[14] = 001_00101100000000000000000
w_carry_translation[14] = 111_10100000000000000000000
{w_sum_translation[14][MSB-1:MSB-2], w_carry_translation[14][MSB-1:MSB-2]} = 01_11 -> q[15] = 0
w[14] = 2 * (w[13] - q[14] * D) = 2 * (
	110_10001100000000000000000 +
	001_11011010000000000000000
) = 2 * 000_01100110000000000000000 = 
000_11001100000000000000000
q_pos = 1000_0010_0100_000
q_neg = 0000_0001_0010_010




// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0111111111100010111011110011 = 134098675
D[WIDTH-1:0] = 0000010000110001000101000011 = 4395331
Q[WIDTH-1:0] = X / D = 30 = 0000000000000000000000011110
REM[WIDTH-1:0] = 134098675 - 4395331 * 30 = 2238745 = 0000001000100010100100011001

CLZ_X = 1
CLZ_D = 5
CLZ_DIFF = CLZ_D - CLZ_X = 4
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 6
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111111111000101110111100110
Divisor[WIDTH-1:0] 		= 1000011000100010100001100000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_000011000100010100001100000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_000110001000101000011000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_111100111011101011110100000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_111001110111010111101000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 010_001000101001000110010000000 >= 0
// 最后一次迭代的商
q[6] = +2
q_pos = 1111_00
q_neg = 0000_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 111100
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 11110
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
0100010001010010001100100000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0100010001010010001100100000 >> 5 = 
0000001000100010100100011001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 0111111111100010111011110011 = 134098675
D[WIDTH-1:0] = 0010000110001000101000011000 = 35162648
Q[WIDTH-1:0] = X / D = 3 = 0000000000000000000000000011
REM[WIDTH-1:0] = 134098675 - 35162648 * 3 = 28610731 = 0001101101001001000010101011

CLZ_X = 1
CLZ_D = 2
CLZ_DIFF = CLZ_D - CLZ_X = 1
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 3
// 最后一次迭代的余数
w[final] = w[3];
w[final] = 011_011010010010000101010110000 >= 0
// 最后一次迭代的商
q[3] = +2
q_pos = 110
q_neg = 000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 110
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 11
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
0110110100100100001010101100
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0110110100100100001010101100 >> 2 = 
0001101101001001000010101011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_111111111000101110111100110
w_sum_translation[0] = w_sum[0] =  001_111111111000101110111100110
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_000000000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_111111110001011101111001100
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_111001110111010111101000000
w_sum_translation[1] = 001_111111110001011101111001100
w_carry_translation[1] = 111_111001110111010111101000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_111111111000101110111100110 +
	110_111100111011101011110100000
) = 2 * 000_111100110100011010110000110 = 
001_111001101000110101100001100
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_111111100010111011110011000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_110011101110101111010000000
w_sum_translation[2] = 001_111111100010111011110011000
w_carry_translation[2] = 001_110011101110101111010000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_01 -> q[3] = +2
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	001_111001101000110101100001100 +
	110_111100111011101011110100000
) = 2 * 001_111001101000110101100001100 = 
011_110011010001101011000011000
q_pos = 110
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_101011110110000110010110000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_101110011011111111000000000
w_sum_translation[3] = 001_101011110110000110010110000
w_carry_translation[3] = 001_101110011011111111000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_01 -> q[4] = +2
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	011_110011010001101011000011000 +
	101_111001110111010111101000000
) = 2 * 001_101101001001000010101011000 = 
011_011010010010000101010110000
q_pos = 1110
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_111000110101011101111100000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
010_101111011101011100000000000
w_sum_translation[4] = 001_111000110101011101111100000
w_carry_translation[4] = 000_101111011101011100000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_00 -> q[5] = +1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	011_011010010010000101010110000 +
	101_111001110111010111101000000
) = 2 * 001_010100001001011100111110000 = 
010_101000010010111001111100000
q_pos = 1110_1
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_010110100111010100010000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_110011110101110111010000000
w_sum_translation[5] = 001_010110100111010100010000000
w_carry_translation[5] = 001_110011110101110111010000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	010_101000010010111001111100000 +
	110_111100111011101011110100000
) = 2 * 001_100101001110100101110000000 = 
011_001010011101001011100000000
q_pos = 1111_00
q_neg = 0000_00

w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_001010011101001011100000000 +
	101_111001110111010111101000000
) = 2 * 001_000100010100100011001000000 = 
010_001000101001000110010000000



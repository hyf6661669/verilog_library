WIDTH = 28
进行R4 SRT迭代时, 需要:
1 + WIDTH + 1 + 2 = 32-bit
来表示"w_sum/w_carry", 其中1-bit是符号位, 1-bit是为了做右移操作的位, 2-bit是初始化的时候要将Dividend右移2位的操作

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110100001110011100100011 = 13690659
D[WIDTH-1:0] = 0000000001001001110111011100 = 302556
Q[WIDTH-1:0] = X / D = 45 = 0000000000000000000000101101
REM[WIDTH-1:0] = 13690659 - 302556 * 45 = 75639 = 0000000000010010011101110111

CLZ_X = 4
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 5
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (6 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(7 / 2) = 4;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 1101000011100111001000110000
Divisor[WIDTH-1:0] 		= 1001001110111011100000000000

+ D = 000_1001001110111011100000000000000
+2D = 001_0010011101110111000000000000000
- D = 111_0110110001000100100000000000000
-2D = 110_1101100010001001000000000000000

4 * (+ D) = 00010_0100111011101110000000000000000
4 * (+2D) = 00100_1001110111011100000000000000000
4 * (- D) = 11101_1011000100010010000000000000000
4 * (-2D) = 11011_0110001000100100000000000000000

根据D的值, 可得选择常数:
m[-1] = -15 = 111_0001
m[ 0] = - 5 = 111_1011
m[+1] = + 5 = 000_0101
m[+2] = +14 = 000_1110

-m[-1]_reduced_2_5 = 00_11110
-m[ 0]_reduced_3_4 = 000_0101
-m[+1]_reduced_3_4 = 111_1011
-m[+2]_reduced_2_5 = 11_00100

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[4];
w[4] = 4 * w[3] - q[4] * D = 
000_1011100010101010011000000000000 + 
111_0110110001000100100000000000000 = 
000_0010010011101110111000000000000 >= 0
// 最后一次迭代的商
q_pos = 0100_0001
q_neg = 0001_0100
corr(q_pos - q_neg) = 00101101

w[final]_reduced >> CLZ_D = 0010010011101110111000000000 >> 9 = 
0000000000010010011101110111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w_sum[0] = 000_0001101000011100111001000110000
w_carry[0] = 000_0000000000000000000000000000000
w[0] = 000_0001101000011100111001000110000
(4 * w[0])_trunc_3_4 = 000_0110, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
111_0000010000110111000100011000000 -> 000_0000010000110111000100011000000
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
000_1101000010000001000000000000000 -> 111_1101000010000001000000000000000
w[1] = 4 * w[0] - q[1] * D = 
000_0110100001110011100100011000000 + 
111_0110110001000100100000000000000 = 
111_1101010010111000000100011000000
(4 * w[1])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[2] = -1

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_10100 + 00_00000 + 00_11110 = 10_10010
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_1010 + 000_0000 + 000_0101 = 001_1111
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_1010 + 000_0000 + 111_1011 = 001_0101
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_10100 + 00_00000 + 11_00100 = 00_11000

(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_10010 + 01_10110)_reduced_2_4 = 
(00_01000)_reduced_2_4 = 00_0100 >= 0
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (001_1111 + 101_1011)_reduced_3_3 = 
(111_1010)_reduced_3_3 = 111_101 < 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (001_0101 + 101_1011)_reduced_3_3 = 
(111_0000)_reduced_3_3 = 111_000 < 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (00_11000 + 01_10110)_reduced_2_4 = 
(10_01110)_reduced_2_4 = 10_0111 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[2] = -1
q_pos = 0100
q_neg = 0001


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
111_1100000101100011110001100000000 -> 000_1100000101100011110001100000000
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
000_0010010100111000000000000000000 -> 111_0010010100111000000000000000000
w[2] = 4 * w[1] - q[2] * D = 
111_0101001011100000010001100000000 + 
000_1001001110111011100000000000000 = 
111_1110011010011011110001100000000
(4 * w[2])_trunc_3_4 = 111_1001, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0100_00
q_neg = 0001_01

// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_01000 + 01_00001 + 00_11110 = 10_00111
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
000_0100 + 101_0000 + 000_0101 = 101_1001
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
000_0100 + 101_0000 + 111_1011 = 100_1111
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_01000 + 01_00001 + 11_00100 = 00_01101


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (10_00111 + 10_01001)_reduced_2_4 = 
(00_10000)_reduced_2_4 = 00_1000 >= 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (101_1001 + 010_0100)_reduced_3_3 = 
(111_1101)_reduced_3_3 = 111_110 < 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (100_1111 + 010_0100)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (00_01101 + 10_01001)_reduced_2_4 = 
(10_10110)_reduced_2_4 = 10_1011 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0100_00
q_neg = 0001_01


ITER[2]:
w[3] = 4 * w[2] - q[3] * D = 
111_1001101001101111000110000000000 + 
000_1001001110111011100000000000000 = 
000_0010111000101010100110000000000
(4 * w[3])_trunc_3_4 = 000_1011, "belongs to [m[+1], m[+2])" -> q[4] = +1
q_pos = 0100_0001
q_neg = 0001_0100

// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_00010 + 10_01010 + 00_11110 = 11_01010
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
100_0001 + 010_0101 + 000_0101 = 110_1011
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
100_0001 + 010_0101 + 111_1011 = 110_0001
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_00010 + 10_01010 + 11_00100 = 01_10000


(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (11_01010 + 10_01001)_reduced_2_4 = 
(01_10011)_reduced_2_4 = 01_1001 >= 0, don't care.
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (110_1011 + 010_0100)_reduced_3_3 = 
(000_1111)_reduced_3_3 = 000_111 >= 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (110_0001 + 010_0100)_reduced_3_3 = 
(000_0101)_reduced_3_3 = 000_010 >= 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (01_10000 + 10_01001)_reduced_2_4 = 
(11_11001)_reduced_2_4 = 11_1100 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[4] = +1
q_pos = 0100_0001
q_neg = 0001_0100



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1111110000100111111000001100 = 264404492
D[WIDTH-1:0] = 0000000000000000000000001001 = 9
Q[WIDTH-1:0] = X / D = 29378276 = 0001110000000100011011100100
REM[WIDTH-1:0] = 264404492 - 9 * 29378276 = 8 = 0000000000000000000000001000
0111000000010001101110010100
CLZ_X = 0
CLZ_D = 24
CLZ_DIFF = CLZ_D - CLZ_X = 24
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (25 % 2) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(26 / 2) = 13;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111110000100111111000001100
Divisor[WIDTH-1:0] 		= 1001000000000000000000000000

+ D = 000_10010000000000000000000000000
+2D = 001_00100000000000000000000000000
- D = 111_01110000000000000000000000000
-2D = 110_11100000000000000000000000000
~ D = 111_01101111111111111111111111111
~2D = 110_11011111111111111111111111111

4 * (+ D) = 00010_01000000000000000000000000000
4 * (+2D) = 00100_10000000000000000000000000000
4 * (- D) = 11101_11000000000000000000000000000
4 * (-2D) = 11011_10000000000000000000000000000

根据D的值, 可得选择常数:
m[-1] = -15 = 111_0001
m[ 0] = - 5 = 111_1011
m[+1] = + 5 = 000_0101
m[+2] = +14 = 000_1110

-m[-1]_reduced_2_5 = 00_11110
-m[ 0]_reduced_3_4 = 000_0101
-m[+1]_reduced_3_4 = 111_1011
-m[+2]_reduced_2_5 = 11_00100

// ---------------------------------------------------------------------------------------------------------------------------------------
w[13] = 4 * w[12] - q[13] * D = 
000_10000000000000000000000000000 + 
111_01110000000000000000000000000 = 
111_11110000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[13];
w[13] = 4 * w[12] - q[13] * D = 
0_10000000000000000000000000000 + 
1_01110000000000000000000000000 = 
1_11110000000000000000000000000 < 0
// 最后一次迭代的商
q_pos = 1000_0000_0001_0010_0000_0001_01
q_neg = 0001_0000_0000_0000_0100_1000_00
corr(q_pos - q_neg) = 0001110000000100011011100100

(w[final]_reduced + (+D)) >> CLZ_D = 
(1111000000000000000000000000 + 1001000000000000000000000000) >> 24 = 
1000000000000000000000000000 >> 24 = 
0000000000000000000000001000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w_sum[0] = 0_0011111100001001111110000011000
w_carry[0] = 0_00000000000000000000000000000
w[0] = 0_0011111100001001111110000011000
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[+2], +Inf)" -> q[1] = +2
q_pos = 10
q_neg = 00


ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
1_10011100001001111110000011000
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_01000000000000000000000000000
w[1] = 4 * w[0] - q[1] * D = 
0_11111100001001111110000011000 + 
0_11100000000000000000000000000 = 
1_11011100001001111110000011000
(4 * w[1])_trunc_3_4 = 111_0111, "belongs to [m[-1], m[0])" -> q[2] = -1

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_11110 + 00_00000 + 00_11110 = 00_11100
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1111 + 000_0000 + 000_0101 = 100_0100
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1111 + 000_0000 + 111_1011 = 011_1010
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_11110 + 00_00000 + 11_00100 = 11_00010


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (00_11100 + 11_10000)_reduced_2_4 = 
(00_01100)_reduced_2_4 = 00_0110 >= 0
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (100_0100 + 011_1000)_reduced_3_3 = 
(111_1100)_reduced_3_3 = 111_110 < 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (011_1010 + 011_1000)_reduced_3_3 = 
(111_0010)_reduced_3_3 = 111_001 < 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (11_00010 + 11_10000)_reduced_2_4 = 
(10_10010)_reduced_2_4 = 10_1001 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[2] = -1
q_pos = 1000
q_neg = 0001


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
1_11100000100111111000001100000
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_00100000000000000000000000000
w[2] = 4 * w[1] - q[2] * D = 
1_01110000100111111000001100000 + 
0_10010000000000000000000000000 = 
0_00000000100111111000001100000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0



// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_11000 + 00_00000 + 00_11110 = 10_10110
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_1100 + 100_0000 + 000_0101 = 110_0001
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_1100 + 100_0000 + 111_1011 = 101_0111
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_11000 + 00_00000 + 11_00100 = 00_11100


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (10_10110 + 10_01000)_reduced_2_4 = 
(00_11110)_reduced_2_4 = 00_1111 >= 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (110_0001 + 010_0100)_reduced_3_3 = 
(000_0101)_reduced_3_3 = 000_010 >= 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (101_0111 + 010_0100)_reduced_3_3 = 
(111_1011)_reduced_3_3 = 111_101 < 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (00_11100 + 10_01000)_reduced_2_4 = 
(11_00100)_reduced_2_4 = 11_0010 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 1000_00
q_neg = 0001_00


ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
1_00000010011111100000110000000
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
1_00000000000000000000000000000
w[3] = 4 * w[2] - q[3] * D = 
0_00000010011111100000110000000 + 
0_00000000000000000000000000000 = 
0_00000010011111100000110000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0

// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_00001 + 10_00000 + 00_11110 = 00_11111
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_0000 + 010_0000 + 000_0101 = 000_0101
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_0000 + 010_0000 + 111_1011 = 111_1011
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_00001 + 10_00000 + 11_00100 = 11_00101

(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (00_11111 + 00_00000)_reduced_2_4 = 
(00_11111)_reduced_2_4 = 00_1111 >= 0, don't care.
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (000_0101 + 000_0000)_reduced_3_3 = 
(000_0101)_reduced_3_3 = 000_010 >= 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (111_1011 + 000_0000)_reduced_3_3 = 
(111_1011)_reduced_3_3 = 111_101 < 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (11_00101 + 00_00000)_reduced_2_4 = 
(11_00101)_reduced_2_4 = 11_0010 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 1000_0000
q_neg = 0001_0000


ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_00001001111110000011000000000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_00000000000000000000000000000
sum + cry = 0_00001001111110000011000000000
w[4] = 4 * w[3] - q[4] * D = 
0_00001001111110000011000000000 + 
0_00000000000000000000000000000 = 
0_00001001111110000011000000000
(4 * w[4])_trunc_3_4 = 000_0010, "belongs to [m[0], m[+1])" -> q[5] = 0


// From the paper:
temp[4][0] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_00100 + 00_00000 + 00_11110 = 01_00010
temp[4][1] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
000_0010 + 000_0000 + 000_0101 = 000_0111
temp[4][2] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
000_0010 + 000_0000 + 111_1011 = 111_1101
temp[4][3] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_00100 + 00_00000 + 11_00100 = 11_01000


(temp[4][0] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (01_00010 + 00_00000)_reduced_2_4 = 
(01_00010)_reduced_2_4 = 01_0001 >= 0, don't care.
(temp[4][1] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (000_0111 + 000_0000)_reduced_3_3 = 
(000_0111)_reduced_3_3 = 000_011 >= 0
(temp[4][2] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (111_1101 + 000_0000)_reduced_3_3 = 
(111_1101)_reduced_3_3 = 111_110 < 0
(temp[4][3] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (11_01000 + 00_00000)_reduced_2_4 = 
(11_01000)_reduced_2_4 = 11_0100 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 1000_0000_00
q_neg = 0001_0000_00


ITER[4]:
w_sum[5] = csa_sum(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
1_00100111111000001100000000000
w_carry[5] = csa_carry(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
1_00000000000000000000000000000
w[5] = 4 * w[4] - q[5] * D = 
0_00100111111000001100000000000 + 
0_00000000000000000000000000000 = 
0_00100111111000001100000000000
(4 * w[5])_trunc_3_4 = 000_1001, "belongs to [m[+1], m[+2])" -> q[6] = +1

// From the paper:
temp[5][0] = ((16 * w_sum[4])_reduced_2_5 + (16 * w_carry[4])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_10011 + 00_00000 + 00_11110 = 01_10001
temp[5][1] = ((16 * w_sum[4])_reduced_3_4 + (16 * w_carry[4])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
000_1001 + 000_0000 + 000_0101 = 000_1110
temp[5][2] = ((16 * w_sum[4])_reduced_3_4 + (16 * w_carry[4])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
000_1001 + 000_0000 + 111_1011 = 000_0100
temp[5][3] = ((16 * w_sum[4])_reduced_2_5 + (16 * w_carry[4])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_10011 + 00_00000 + 11_00100 = 11_10111

(temp[5][0] + (-4 * q[5] * D)_reduced_2_5)_reduced_2_4 = (01_10001 + 00_00000)_reduced_2_4 = 
(01_10001)_reduced_2_4 = 01_1000 >= 0, don't care.
(temp[5][1] + (-4 * q[5] * D)_reduced_3_4)_reduced_3_3 = (000_1110 + 000_0000)_reduced_3_3 = 
(000_1110)_reduced_3_3 = 000_111 >= 0
(temp[5][2] + (-4 * q[5] * D)_reduced_3_4)_reduced_3_3 = (000_0100 + 000_0000)_reduced_3_3 = 
(000_0100)_reduced_3_3 = 000_010 >= 0
(temp[5][3] + (-4 * q[5] * D)_reduced_2_5)_reduced_2_4 = (11_10111 + 00_00000)_reduced_2_4 = 
(11_10111)_reduced_2_4 = 11_1011 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[6] = +1
q_pos = 1000_0000_0001
q_neg = 0001_0000_0000


ITER[5]:
w_sum[6] = csa_sum(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
1_11101111100000110000000000000
w_carry[6] = csa_carry(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
0_00100000000000000000000000000
w[6] = 4 * w[5] - q[6] * D = 
0_10011111100000110000000000000 + 
1_01110000000000000000000000000 = 
0_00001111100000110000000000000
(4 * w[6])_trunc_3_4 = 000_0011, "belongs to [m[0], m[+1])" -> q[7] = 0

// From the paper:
temp[6][0] = ((16 * w_sum[5])_reduced_2_5 + (16 * w_carry[5])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_01111 + 00_00000 + 00_11110 = 11_01101
temp[6][1] = ((16 * w_sum[5])_reduced_3_4 + (16 * w_carry[5])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
010_0111 + 000_0000 + 000_0101 = 010_1100
temp[6][2] = ((16 * w_sum[5])_reduced_3_4 + (16 * w_carry[5])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
010_0111 + 000_0000 + 111_1011 = 010_0010
temp[6][3] = ((16 * w_sum[5])_reduced_2_5 + (16 * w_carry[5])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_01111 + 00_00000 + 11_00100 = 01_10011


(temp[6][0] + (-4 * q[6] * D)_reduced_2_5)_reduced_2_4 = (11_01101 + 01_11000)_reduced_2_4 = 
(01_00101)_reduced_2_4 = 01_0010 >= 0, don't care.
(temp[6][1] + (-4 * q[6] * D)_reduced_3_4)_reduced_3_3 = (010_1100 + 101_1100)_reduced_3_3 = 
(000_1000)_reduced_3_3 = 000_100 >= 0
(temp[6][2] + (-4 * q[6] * D)_reduced_3_4)_reduced_3_3 = (010_0010 + 101_1100)_reduced_3_3 = 
(111_1110)_reduced_3_3 = 111_111 < 0
(temp[6][3] + (-4 * q[6] * D)_reduced_2_5)_reduced_2_4 = (01_10011 + 01_11000)_reduced_2_4 = 
(11_01011)_reduced_2_4 = 11_0101 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 1000_0000_0001_00
q_neg = 0001_0000_0000_00


ITER[6]:
w_sum[7] = csa_sum(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
1_00111110000011000000000000000
w_carry[7] = csa_carry(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
1_00000000000000000000000000000
w[7] = 4 * w[6] - q[7] * D = 
0_00111110000011000000000000000 + 
0_00000000000000000000000000000 = 
0_00111110000011000000000000000
(4 * w[7])_trunc_3_4 = 000_1111, "belongs to [m[+2], +Inf)" -> q[8] = +2

// From the paper:
temp[7][0] = ((16 * w_sum[6])_reduced_2_5 + (16 * w_carry[6])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_11111 + 10_00000 + 00_11110 = 01_11101
temp[7][1] = ((16 * w_sum[6])_reduced_3_4 + (16 * w_carry[6])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_1111 + 010_0000 + 000_0101 = 001_0100
temp[7][2] = ((16 * w_sum[6])_reduced_3_4 + (16 * w_carry[6])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_1111 + 010_0000 + 111_1011 = 000_1010
temp[7][3] = ((16 * w_sum[6])_reduced_2_5 + (16 * w_carry[6])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_11111 + 10_00000 + 11_00100 = 00_00011


(temp[7][0] + (-4 * q[7] * D)_reduced_2_5)_reduced_2_4 = (01_11101 + 00_00000)_reduced_2_4 = 
(01_11101)_reduced_2_4 = 01_1110 >= 0, don't care.
(temp[7][1] + (-4 * q[7] * D)_reduced_3_4)_reduced_3_3 = (001_0100 + 000_0000)_reduced_3_3 = 
(001_0100)_reduced_3_3 = 001_010 >= 0
(temp[7][2] + (-4 * q[7] * D)_reduced_3_4)_reduced_3_3 = (000_1010 + 000_0000)_reduced_3_3 = 
(000_1010)_reduced_3_3 = 000_101 >= 0
(temp[7][3] + (-4 * q[7] * D)_reduced_2_5)_reduced_2_4 = (00_00011 + 00_00000)_reduced_2_4 = 
(00_00011)_reduced_2_4 = 00_0001 >= 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 1000_0000_0001_0010
q_neg = 0001_0000_0000_0000


ITER[7]:
w_sum[8] = csa_sum(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
0_00011000001100000000000000000
w_carry[8] = csa_carry(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
1_11000000000000000000000000000
w[8] = 4 * w[7] - q[8] * D = 
0_11111000001100000000000000000 + 
0_11100000000000000000000000000 = 
1_11011000001100000000000000000
(4 * w[8])_trunc_3_4 = 111_0110, "belongs to [m[-1], m[0])" -> q[9] = -1

// From the paper:
temp[8][0] = ((16 * w_sum[7])_reduced_2_5 + (16 * w_carry[7])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_11100 + 00_00000 + 00_11110 = 00_11010
temp[8][1] = ((16 * w_sum[7])_reduced_3_4 + (16 * w_carry[7])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1110 + 000_0000 + 000_0101 = 100_0011
temp[8][2] = ((16 * w_sum[7])_reduced_3_4 + (16 * w_carry[7])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1110 + 000_0000 + 111_1011 = 011_1001
temp[8][3] = ((16 * w_sum[7])_reduced_2_5 + (16 * w_carry[7])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_11100 + 00_00000 + 11_00100 = 11_00000


(temp[8][0] + (-4 * q[8] * D)_reduced_2_5)_reduced_2_4 = (00_11010 + 11_10000)_reduced_2_4 = 
(00_01010)_reduced_2_4 = 00_0101 >= 0
(temp[8][1] + (-4 * q[8] * D)_reduced_3_4)_reduced_3_3 = (100_0011 + 011_1000)_reduced_3_3 = 
(111_1011)_reduced_3_3 = 111_101 < 0
(temp[8][2] + (-4 * q[8] * D)_reduced_3_4)_reduced_3_3 = (011_1001 + 011_1000)_reduced_3_3 = 
(111_0001)_reduced_3_3 = 111_000 < 0
(temp[8][3] + (-4 * q[8] * D)_reduced_2_5)_reduced_2_4 = (11_00000 + 11_10000)_reduced_2_4 = 
(10_10000)_reduced_2_4 = 10_1000 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[9] = -1
q_pos = 1000_0000_0001_0010_00
q_neg = 0001_0000_0000_0000_01

ITER[8]:
w_sum[9] = csa_sum(4 * w_sum[8], 4 * w_carry[8], -q[9] * D) = 
1_11110000110000000000000000000
w_carry[9] = csa_carry(4 * w_sum[8], 4 * w_carry[8], -q[9] * D) = 
0_00000000000000000000000000000
w[9] = 4 * w[8] - q[9] * D = 
1_01100000110000000000000000000 + 
0_10010000000000000000000000000 = 
1_11110000110000000000000000000
(4 * w[9])_trunc_3_4 = 111_1100, "belongs to [m[0], m[+1])" -> q[10] = 0

// From the paper:
temp[9][0] = ((16 * w_sum[8])_reduced_2_5 + (16 * w_carry[8])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_10000 + 00_00000 + 00_11110 = 10_01110
temp[9][1] = ((16 * w_sum[8])_reduced_3_4 + (16 * w_carry[8])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_1000 + 100_0000 + 000_0101 = 101_1101
temp[9][2] = ((16 * w_sum[8])_reduced_3_4 + (16 * w_carry[8])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_1000 + 100_0000 + 111_1011 = 101_0011
temp[9][3] = ((16 * w_sum[8])_reduced_2_5 + (16 * w_carry[8])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_10000 + 00_00000 + 11_00100 = 00_10100


(temp[9][0] + (-4 * q[9] * D)_reduced_2_5)_reduced_2_4 = (10_01110 + 10_01000)_reduced_2_4 = 
(00_10110)_reduced_2_4 = 00_1011 >= 0, don't care.
(temp[9][1] + (-4 * q[9] * D)_reduced_3_4)_reduced_3_3 = (101_1101 + 010_0100)_reduced_3_3 = 
(000_0001)_reduced_3_3 = 000_000 >= 0
(temp[9][2] + (-4 * q[9] * D)_reduced_3_4)_reduced_3_3 = (101_0011 + 010_0100)_reduced_3_3 = 
(111_0111)_reduced_3_3 = 111_011 < 0
(temp[9][3] + (-4 * q[9] * D)_reduced_2_5)_reduced_2_4 = (00_10100 + 10_01000)_reduced_2_4 = 
(10_11100)_reduced_2_4 = 10_1110 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 1000_0000_0001_0010_0000
q_neg = 0001_0000_0000_0000_0100


ITER[9]:
w_sum[10] = csa_sum(4 * w_sum[9], 4 * w_carry[9], -q[10] * D) = 
1_11000011000000000000000000000
w_carry[10] = csa_carry(4 * w_sum[9], 4 * w_carry[9], -q[10] * D) = 
0_00000000000000000000000000000
w[10] = 4 * w[9] - q[10] * D = 
1_11000011000000000000000000000 + 
0_00000000000000000000000000000 = 
1_11000011000000000000000000000
(4 * w[10])_trunc_3_4 = 111_0000, "belongs to (-Inf, m[-1])" -> q[11] = -2

// From the paper:
temp[10][0] = ((16 * w_sum[9])_reduced_2_5 + (16 * w_carry[9])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_00001 + 00_00000 + 00_11110 = 11_11111
temp[10][1] = ((16 * w_sum[9])_reduced_3_4 + (16 * w_carry[9])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
111_0000 + 000_0000 + 000_0101 = 111_0101
temp[10][2] = ((16 * w_sum[9])_reduced_3_4 + (16 * w_carry[9])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
111_0000 + 000_0000 + 111_1011 = 110_1011
temp[10][3] = ((16 * w_sum[9])_reduced_2_5 + (16 * w_carry[9])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_00001 + 00_00000 + 11_00100 = 10_00101


(temp[10][0] + (-4 * q[10] * D)_reduced_2_5)_reduced_2_4 = (11_11111 + 00_00000)_reduced_2_4 = 
(11_11111)_reduced_2_4 = 11_1111 < 0
(temp[10][1] + (-4 * q[10] * D)_reduced_3_4)_reduced_3_3 = (111_0101 + 000_0000)_reduced_3_3 = 
(111_0101)_reduced_3_3 = 111_010 < 0
(temp[10][2] + (-4 * q[10] * D)_reduced_3_4)_reduced_3_3 = (110_1011 + 000_0000)_reduced_3_3 = 
(110_1011)_reduced_3_3 = 110_101 < 0
(temp[10][3] + (-4 * q[10] * D)_reduced_2_5)_reduced_2_4 = (10_00101 + 00_00000)_reduced_2_4 = 
(10_00101)_reduced_2_4 = 10_0010 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to (-Inf, m[-1])" -> q[11] = -2
q_pos = 1000_0000_0001_0010_0000_00
q_neg = 0001_0000_0000_0000_0100_10


ITER[10]:
w_sum[11] = csa_sum(4 * w_sum[10], 4 * w_carry[10], -q[11] * D) = 
0_00101100000000000000000000000
w_carry[11] = csa_carry(4 * w_sum[10], 4 * w_carry[10], -q[11] * D) = 
0_00000000000000000000000000000
w[11] = 4 * w[10] - q[11] * D = 
1_00001100000000000000000000000 + 
1_00100000000000000000000000000 = 
0_00101100000000000000000000000
(4 * w[11])_trunc_3_4 = 000_1011, "belongs to [m[+1], m[+2])" -> q[12] = +1

// From the paper:
temp[11][0] = ((16 * w_sum[10])_reduced_2_5 + (16 * w_carry[10])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_00110 + 00_00000 + 00_11110 = 01_00100
temp[11][1] = ((16 * w_sum[10])_reduced_3_4 + (16 * w_carry[10])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
100_0011 + 000_0000 + 000_0101 = 100_1000
temp[11][2] = ((16 * w_sum[10])_reduced_3_4 + (16 * w_carry[10])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
100_0011 + 000_0000 + 111_1011 = 011_1110
temp[11][3] = ((16 * w_sum[10])_reduced_2_5 + (16 * w_carry[10])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_00110 + 00_00000 + 11_00100 = 11_01010


(temp[11][0] + (-4 * q[11] * D)_reduced_2_5)_reduced_2_4 = (01_00100 + 00_10000)_reduced_2_4 = 
(01_10100)_reduced_2_4 = 01_1010 >= 0, don't care.
(temp[11][1] + (-4 * q[11] * D)_reduced_3_4)_reduced_3_3 = (100_1000 + 100_1000)_reduced_3_3 = 
(001_0000)_reduced_3_3 = 001_000 >= 0
(temp[11][2] + (-4 * q[11] * D)_reduced_3_4)_reduced_3_3 = (011_1110 + 100_1000)_reduced_3_3 = 
(000_0110)_reduced_3_3 = 000_011 >= 0
(temp[11][3] + (-4 * q[11] * D)_reduced_2_5)_reduced_2_4 = (11_01010 + 00_10000)_reduced_2_4 = 
(11_11010)_reduced_2_4 = 11_1101 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[12] = +1
q_pos = 1000_0000_0001_0010_0000_0001
q_neg = 0001_0000_0000_0000_0100_1000


ITER[11]:
w_sum[12] = csa_sum(4 * w_sum[11], 4 * w_carry[11], -q[12] * D) = 
1_11000000000000000000000000000
w_carry[12] = csa_carry(4 * w_sum[11], 4 * w_carry[11], -q[12] * D) = 
0_01100000000000000000000000000
w[12] = 4 * w[11] - q[12] * D = 
0_10110000000000000000000000000 + 
1_01110000000000000000000000000 = 
0_00100000000000000000000000000
(4 * w[12])_trunc_3_4 = 000_1011, "belongs to [m[+1], m[+2])" -> q[13] = +1

// From the paper:
temp[12][0] = ((16 * w_sum[11])_reduced_2_5 + (16 * w_carry[11])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_11000 + 00_00000 + 00_11110 = 11_10110
temp[12][1] = ((16 * w_sum[11])_reduced_3_4 + (16 * w_carry[11])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
010_1100 + 000_0000 + 000_0101 = 011_0001
temp[12][2] = ((16 * w_sum[11])_reduced_3_4 + (16 * w_carry[11])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
010_1100 + 000_0000 + 111_1011 = 010_0111
temp[12][3] = ((16 * w_sum[11])_reduced_2_5 + (16 * w_carry[11])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_11000 + 00_00000 + 11_00100 = 01_11100


(temp[12][0] + (-4 * q[12] * D)_reduced_2_5)_reduced_2_4 = (11_10110 + 01_11000)_reduced_2_4 = 
(01_01110)_reduced_2_4 = 01_0111 >= 0, don't care.
(temp[12][1] + (-4 * q[12] * D)_reduced_3_4)_reduced_3_3 = (011_0001 + 101_1100)_reduced_3_3 = 
(000_1101)_reduced_3_3 = 000_110 >= 0
(temp[12][2] + (-4 * q[12] * D)_reduced_3_4)_reduced_3_3 = (010_0111 + 101_1100)_reduced_3_3 = 
(000_0011)_reduced_3_3 = 000_001 >= 0
(temp[12][3] + (-4 * q[12] * D)_reduced_2_5)_reduced_2_4 = (01_11100 + 01_11000)_reduced_2_4 = 
(11_10100)_reduced_2_4 = 11_1010 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[13] = +1
q_pos = 1000_0000_0001_0010_0000_0001_01
q_neg = 0001_0000_0000_0000_0100_1000_00






接"test_1.sv".

最后试了N多个例子, 发现如果"q[final] = -1/+1", 则会导致无法求出正确的余数, 所以还是简单粗暴一点, 要求"WIDTH-bit"整数除法的商和余数时, 只做"(WIDTH + 1)"
次迭代.
// ---------------------------------------------------------------------------------------------------------------------------------------
先考虑无符号整数除法，根据论文对其算法的属性的描述，以及从下面的例子可以得到如下结论:
Q[final]: 最后一次迭代得到的商的非冗余形式.
w[final] = w_sum[final] + w_carry[final];
W[final] = w[final] / 2;
quotient: 商的绝对值.
remainder: 余数的绝对值.
有以下几种情况:
1. W[final]属于区间"[+ D, +2D)" -> quotient = Q[final] + 1, remainder = (W[final] -  D) >> CLZ_D;
2. W[final]属于区间"[+ 0, + D)" -> quotient = Q[final] + 0, remainder = (W[final] +  0) >> CLZ_D;
3. W[final]属于区间"[- D, - 0)" -> quotient = Q[final] - 1, remainder = (W[final] +  D) >> CLZ_D;
4. W[final]属于区间"[-2D, - D)" -> quotient = Q[final] - 2, remainder = (W[final] + 2D) >> CLZ_D;
总的来说, 大致需要7个全加计算:
fa[0] = w_sum + w_carry;
fa[1] = fa[0] + (-D);
fa[2] = fa[0] + D;
fa[3] = fa[0] + 2D;
fa[4] = Q[final] + 1;
fa[5] = Q[final] - 1;
fa[6] = Q[final] - 2;


Q[0] = 1: Q - 1'b1 = {Q[WIDTH-1:1] - 1'b0, 1'b0} = {Q[WIDTH-1:1], ~Q[0]};
Q[0] = 0: Q - 1'b1 = {Q[WIDTH-1:1] - 1'b1, 1'b1} = {Q[WIDTH-1:1] - 1'b1, ~Q[0]};
Q - 2 = Q - 2'b10 = {Q[WIDTH-1:1] - 1'b1, Q[0]};

由上述等式可知, 在计算"fa[6], fa[5]"时, 可以使用"1个full adder + 1个MUX"来代替"2个full adder", 可能会有某种收益.

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
对于有符号数除法来说, 当余数为负数时(余数和被除数"Dividend"同号, 在前处理过程中就知道余数是否应该为负数), 有类似的结论.
Q[final]: 最后一次迭代得到的商的非冗余形式, 绝对值.
w[final] = (-w_sum_translation[final]) + (-w_carry_translation[final]) =
~w_sum_translation[final] + ~w_carry_translation[final] + 2'b10;
W[final] = w[final] / 2;
quotient: 修正后的商, 绝对值.
remainder: 修正后的余数, 有符号数.
1. W[final]属于区间"(-2D, - D]" -> quotient = Q[final] + 1, remainder = (W[final] +  D) >> CLZ_D;
2. W[final]属于区间"(- D, - 0]" -> quotient = Q[final] + 0, remainder = (W[final] +  0) >> CLZ_D;
3. W[final]属于区间"(+ 0, + D]" -> quotient = Q[final] - 1, remainder = (W[final] -  D) >> CLZ_D;
4. W[final]属于区间"(+ D, +2D]" -> quotient = Q[final] - 2, remainder = (W[final] - 2D) >> CLZ_D;
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
post_process最主要的目标是:
1. 余数为非正数 -> 计算出属于区间"(-D, -0]"的"remainder".
2. 余数为非负数 -> 计算出属于区间"[+0, +D)"的"remainder".
因此"Q[final] + 1, Q[final] - 1, Q[final] - 2"都属于"Speculative(预测性的)"计算.为了减少FA的数量，可以在后处理中先算出修正后的remainder, 然后根据修正操作时
使用到的系数(+2/-2, +1/-1, 0)计算出最终的quotient. 于是可将后处理分为2步:
1. 并行计算"W[fianl], W[final] + D, W[final] + (-D), (W[final] + 2D)(余数为非负数)/(W[final] - 2D)(余数为非正数)".
2. 对修正后的"W[final]"进行右移操作得到正确的余数"remainder", 根据步骤1中的系数计算出正确的商quotient.
大致可将步骤1和步骤2分别放在2个周期里完成.

综上所述, 每一步主要需要的运算器包括:
1. pre_process.
2个"WIDTH-bit"的FA: 计算被除数和除数的绝对值.
2个lzc: 计算被除数和除数的绝对值的前导0个数.
2个left_shifter: 根据LZC对被除数和除数进行左移.

2. srt_iter, 以"4个Radix-2叠加起来形成Radix-16"为例.
1个"(WIDTH - 4)-bit"的FA: 计算上次大迭代得到的商数字的非冗余形式.
2个"4-bit"的FA: 计算本次大迭代前3次小迭代得到的商数字的非冗余形式.

3. post_process.
4个"(WIDTH + 2)-bit"的FA: 确定"W[final] = w[final] / 2"属于哪个区间.
1个"WIDTH-bit"的FA: 计算quotient, post_process_0先算remainder_pre, post_process_1再计算quotient, 所以不需要为计算quotient分配独立的FA.
1个right_shifter: 计算remainder, 可以和pre_process中的left_shifter复用.

综上所述, 一共需要:
4个"(WIDTH + 2)-bit"的FA.
2个lzc.
2个left_shifter.
若干个CSA, MUX.....

// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000010000000110000 = 8240
Q[WIDTH-1:0] = X / D = 87 = 000000000000000001010111
REM[WIDTH-1:0] = 717047 - 8240 * 87 = 167 = 000000000000000010100111

CLZ_X = 4
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 6
迭代次数:
iter_num = CLZ_DIFF + 1 = 7
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101011110000111101110000
Divisor[WIDTH-1:0] 		= 100000001100000000000000

+ D[(WIDTH + 2)-1:0] = 001_00000001100000000000000
+2D[(WIDTH + 2)-1:0] = 010_00000011000000000000000
- D[(WIDTH + 2)-1:0] = 110_11111110100000000000000
-2D[(WIDTH + 2)-1:0] = 101_11111101000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[7] = 010_00001101011100000000000 > 0
w[final] / 2 + (-D) = 
001_00000110101110000000000 + 110_11111110100000000000000 = 
000_00000101001110000000000 > 0 -> (w[final] / 2) "belongs to [+D, +2D)".
// 最后一次迭代的商
q_pos = 1010_110
q_neg = 0000_000

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 1010110;
(w[final] / 2) "belongs to [+ D, +2D)" -> quotient_correction_coefficient = 1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 1010111;

(w[final] / 2) "belongs to [+ D, +2D)" -> remainder_correction_coefficient = 1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
000000101001110000000000 >> 10 = 
000000000000000010100111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 余数是负数
REM[WIDTH-1:0] = -167 = 111111111111111101011001

w_sum_translation[final] = 000_00111001011100000000000
w_carry_translation[final] = 001_11010100000000000000000
~w_sum_translation[final] = 111_11000110100011111111111
~w_carry_translation[final] = 110_00101011111111111111111

w[final] = ~w_sum_translation[final] + ~w_carry_translation[final] + 2'b10 = 101_11110010100100000000000 < 0
(w[final] / 2) + D = 110_11111001010010000000000 + 001_00000001100000000000000 = 
111_11111010110010000000000 < 0 -> (w[final] / 2) "belongs to (-2D, -D]".

remainder_calculated[WIDTH-1:0] = ((w[final] / 2) + D) >> CLZ_D = 
(110_11111001010010000000000 + 001_00000001100000000000000) >> 10 = 
111_11111010110010000000000 >> 10 = 
111111111111111101011001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000100000001100000000 = 131840
Q[WIDTH-1:0] = X / D = 5 = 000000000000000000000101
REM[WIDTH-1:0] = 717047 - 131840 * 5 = 57847 = 000000001110000111110111

CLZ_X = 4
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 2
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 4
q[3] = 0
q[4] = +1
q_pos = 1001
q_neg = 0000
q_pos - q_neg = 1001
w[4] = 011_11000110111011100000000 >= 0
w[4] / 2 = 001_11100011011101110000000
001_11100011011101110000000 + (-D) = 
001_11100011011101110000000 + 110_11111110100000000000000 = 
000_11100001111101110000000

011100001111101110000000 >> (CLZ_D + 1) = 
000000001110000111110111
// ---------------------------------------------------------------------------------------------------------------------------------------




初始化:
w[0][(WIDTH + 2)-1:0] = 001_01011110000111101110000
w_sum_translation[0] = w_sum[0] = 001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_10111100001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11111101000000000000000
w_sum_translation[1] = 000_10111100001111011100000
w_carry_translation[1] = 111_11111101000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01011110000111101110000 +
	110_11111110100000000000000
) = 2 * 000_01011100100111101110000 = 
000_10111001001111011100000
q_pos = 10
q_neg = 00


w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_01111000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11111010000000000000000
w_sum_translation[2] = 001_01111000011110111000000
w_carry_translation[2] = 111_11111010000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_10111001001111011100000 +
	000_00000000000000000000000
) = 2 * 000_10111001001111011100000 = 
001_01110010011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_11110000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_11110100000000000000000
w_sum_translation[3] = 000_11110000111101110000000
w_carry_translation[3] = 001_11110100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_01 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_01110010011110111000000 +
	000_00000000000000000000000
) = 2 * 001_01110010011110111000000 = 
010_11100100111101110000000
q_pos = 1001
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_11110100111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11010010000000000000000
w_sum_translation[4] = 001_11110100111011100000000
w_carry_translation[4] = 001_11010010000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[5] = +2
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	010_11100100111101110000000 +
	110_11111110100000000000000
) = 2 * 001_11100011011101110000000 = 
011_11000110111011100000000
q_pos = 1010_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_10110111110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11010000000000000000000
w_sum_translation[5] = 001_10110111110111000000000
w_carry_translation[5] = 001_11010000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	011_11000110111011100000000 +
	101_11111101000000000000000
) = 2 * 001_11000011111011100000000 = 
011_10000111110111000000000
q_pos = 1010_10
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_00110101101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_11010100000000000000000
w_sum_translation[6] = 001_00110101101110000000000
w_carry_translation[6] = 001_11010100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_01 -> q[7] = +2
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_10000111110111000000000 +
	101_11111101000000000000000
) = 2 * 001_10000100110111000000000 = 
011_00001001101110000000000
q_pos = 1010_110
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_00111001011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_11010100000000000000000
w_sum_translation[7] = 000_00111001011100000000000
w_carry_translation[7] = 001_11010100000000000000000
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	011_00001001101110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000110101110000000000 = 
010_00001101011100000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000000010101011 = 171
Q[WIDTH-1:0] = X / D = 4193 = 000000000001000001100001
REM[WIDTH-1:0] = 717047 - 171 * 4193 = 44 = 000000000000000000101100

CLZ_X = 4
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 12
迭代次数:
iter_num = CLZ_DIFF + 1 = 13
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101011110000111101110000
Divisor[WIDTH-1:0] 		= 101010110000000000000000

+ D[(WIDTH + 2)-1:0] = 001_01010110000000000000000
+2D[(WIDTH + 2)-1:0] = 010_10101100000000000000000
- D[(WIDTH + 2)-1:0] = 110_10101010000000000000000
-2D[(WIDTH + 2)-1:0] = 101_01010100000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[13] = 000_10110000000000000000000 >= 0
(w[final] / 2) + (-D) = 000_01011000000000000000000 + 110_10101010000000000000000 = 
11100000010000000000000000 < 0 -> (w[final] / 2) "belongs to [+0, +D)";
001011000000000000000000
// 最后一次迭代的商
q_pos = 1000_0100_0000_0
q_neg = 0000_0000_1111_1

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 0001000001100001;
(w[final] / 2) "belongs to [+0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 0001000001100001;

(w[final] / 2) "belongs to [+0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
001011000000000000000000 >> 16 = 
000000000000000000101100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 余数是负数
REM[WIDTH-1:0] = -44 = 111111111111111111010100

w_sum_translation[final] = 001_01001000000000000000000
w_carry_translation[final] = 111_01101000000000000000000
~w_sum_translation[final] = 110_10110111111111111111111
~w_carry_translation[final] = 000_10010111111111111111111

w[final] = ~w_sum_translation[final] + ~w_carry_translation[final] + 2'b10 = 111_01010000000000000000000 < 0
(w[final] / 2) + D = 111_10101000000000000000000 + 001_01010110000000000000000 = 
000_11111110000000000000000 >= 0 -> (w[final] / 2) "belongs to (-D, -0]".

remainder_calculated[WIDTH-1:0] = ((w[final] / 2) + 0) >> CLZ_D = 
110101000000000000000000 >> 16 = 
111111111111111111010100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000001010101100000000 = 43776
Q[WIDTH-1:0] = X / D = 16 = 000000000000000000010000
REM[WIDTH-1:0] = 717047 - 43776 * 16 = 16631 = 000000000100000011110111

CLZ_X = 4
CLZ_D = 8
CLZ_DIFF = CLZ_D - CLZ_X = 4
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 6
q[5] = 0
q[6] = +1
q_pos = 1000_01
q_neg = 0000_00
q_pos - q_neg = 100001
w[6] = 111_01011011101110000000000
w[6] / 2 = 111_10101101110111000000000
111_10101101110111000000000 + (D) = 
111_10101101110111000000000 + 001_01010110000000000000000 = 
001_00000011110111000000000

100000011110111000000000 >> (CLZ_D + 1) = 
000000000100000011110111

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000001010101100000 = 5472
Q[WIDTH-1:0] = X / D = 131 = 000000000000000010000011
REM[WIDTH-1:0] = 717047 - 5472 * 131 = 215 = 000000000000000011010111

CLZ_X = 4
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 7
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 9
q[8] = 0
q[9] = -1
q_pos = 1000_0100_0
q_neg = 0000_0000_1
q_pos - q_neg = 000100000111
w[9] = 101_10001001110000000000000 < 0
w[9] / 2 = 110_11000100111000000000000
110_11000100111000000000000 + (D) = 
110_11000100111000000000000 + 001_01010110000000000000000 = 
000_00011010111000000000000

000011010111000000000000 >> (CLZ_D + 1) = 
000000000000000011010111

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000000101010110 = 342
Q[WIDTH-1:0] = X / D = 2096 = 000000000000100000110000
REM[WIDTH-1:0] = 717047 - 342 * 2096 = 215 = 000000000000000011010111

CLZ_X = 4
CLZ_D = 15
CLZ_DIFF = CLZ_D - CLZ_X = 11
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 13
q[12] = -1
q[13] = -1
q_pos = 1000_0100_0000_0
q_neg = 0000_0000_1111_1
q_pos - q_neg = 0001000001100001

w[13] = 000_10110000000000000000000 >= 0
w[13] / 2 = 000_01011000000000000000000
000_01011000000000000000000 + (D) = 
000_01011000000000000000000 + 001_01010110000000000000000 = 
110101110000000000000000

110101110000000000000000 >> (CLZ_D + 1) = 
000000000000000011010111

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000001010101100 = 684
Q[WIDTH-1:0] = X / D = 1048 = 000000000000010000011000
REM[WIDTH-1:0] = 717047 - 684 * 1048 = 215 = 000000000000000011010111

CLZ_X = 4
CLZ_D = 14
CLZ_DIFF = CLZ_D - CLZ_X = 10
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 12
q[11] = -1
q[12] = -1
q_pos = 1000_0100_0000
q_neg = 0000_0000_1111
q_pos - q_neg = 100000110001
w[12] = 111_00000010000000000000000 < 0
w[12] / 2 = 111_10000001000000000000000
111_10000001000000000000000 + (D) = 
111_10000001000000000000000 + 001_01010110000000000000000 = 
000_11010111000000000000000

011010111000000000000000 >> (CLZ_D + 1) = 
000000000000000011010111

// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 2)-1:0] =  001_01011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
111_11101000001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_00101000000000000000000
w_sum_translation[1] = 111_11101000001111011100000
w_carry_translation[1] = 000_00101000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_00 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01011110000111101110000 +
	110_10101010000000000000000
) = 2 * 000_00001000000111101110000 = 
000_00010000001111011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11010000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_01010000000000000000000
w_sum_translation[2] = 111_11010000011110111000000
w_carry_translation[2] = 000_01010000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 11_00 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_00010000001111011100000 +
	000_00000000000000000000000
) = 2 * 000_00010000001111011100000 = 
000_00100000011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_10100000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_10100000000000000000000
w_sum_translation[3] = 111_10100000111101110000000
w_carry_translation[3] = 000_10100000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_00 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00100000011110111000000 +
	000_00000000000000000000000
) = 2 * 000_00100000011110111000000 = 
000_01000000111101110000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_01000001111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_01000000000000000000000
w_sum_translation[4] = 111_01000001111011100000000
w_carry_translation[4] = 001_01000000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_01 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_01000000111101110000000 +
	000_00000000000000000000000
) = 2 * 000_01000000111101110000000 = 
000_10000001111011100000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_10000011110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
010_10000000000000000000000
w_sum_translation[5] = 000_10000011110111000000000
w_carry_translation[5] = 000_10000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_00 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_10000001111011100000000 +
	000_00000000000000000000000
) = 2 * 000_10000001111011100000000 = 
001_00000011110111000000000
q_pos = 1000_01
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_01010011101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
110_00001000000000000000000
w_sum_translation[6] = 001_01010011101110000000000
w_carry_translation[6] = 110_00001000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	001_00000011110111000000000 +
	110_10101010000000000000000
) = 2 * 111_10101101110111000000000 = 
111_01011011101110000000000
q_pos = 1000_010
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_10100111011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
100_00010000000000000000000
w_sum_translation[7] = 000_10100111011100000000000
w_carry_translation[7] = 110_00010000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_10 -> q[8] = 0
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	111_01011011101110000000000 +
	000_00000000000000000000000
) = 2 * 111_01011011101110000000000 = 
110_10110111011100000000000
q_pos = 1000_0100
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
001_01001110111000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
100_00100000000000000000000
w_sum_translation[8] = 111_01001110111000000000000
w_carry_translation[8] = 110_00100000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 11_10 -> q[9] = -1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	110_10110111011100000000000 +
	000_00000000000000000000000
) = 2 * 110_10110111011100000000000 = 
101_01101110111000000000000
q_pos = 1000_0100_0
q_neg = 0000_0000_1

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
100_01110001110000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
001_00011000000000000000000
w_sum_translation[9] = 110_01110001110000000000000
w_carry_translation[9] = 111_00011000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_11 -> q[10] = -1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	101_01101110111000000000000 +
	001_01010110000000000000000
) = 2 * 110_11000100111000000000000 = 
101_10001001110000000000000
q_pos = 1000_0100_00
q_neg = 0000_0000_11

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
100_01111111100000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_01000000000000000000000
w_sum_translation[10] = 110_01111111100000000000000
w_carry_translation[10] = 111_01000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 10_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	101_10001001110000000000000 +
	001_01010110000000000000000
) = 2 * 110_11011111110000000000000 = 
101_10111111100000000000000
q_pos = 1000_0100_000
q_neg = 0000_0000_111

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_11010011000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
001_01011000000000000000000
w_sum_translation[11] = 110_11010011000000000000000
w_carry_translation[11] = 111_01011000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_11 -> q[12] = -1
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	101_10111111100000000000000 +
	001_01010110000000000000000
) = 2 * 111_00010101100000000000000 = 
110_00101011000000000000000
q_pos = 1000_0100_0000
q_neg = 0000_0000_1111

w_sum[12] = 2 * csa_sum(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
101_10111010000000000000000
w_carry[12] = 2 * csa_carry(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
001_01001000000000000000000
w_sum_translation[12] = 111_10111010000000000000000
w_carry_translation[12] = 111_01001000000000000000000
{w_sum_translation[12][MSB-1:MSB-2], w_carry_translation[12][MSB-1:MSB-2]} = 11_11 -> q[13] = -1
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	110_00101011000000000000000 +
	001_01010110000000000000000
) = 2 * 111_10000001000000000000000 = 
111_00000010000000000000000
q_pos = 1000_0100_0000_0
q_neg = 0000_0000_1111_1

w_sum[13] = 2 * csa_sum(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
011_01001000000000000000000
w_carry[13] = 2 * csa_carry(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
101_01101000000000000000000
w_sum_translation[13] = 001_01001000000000000000000
w_carry_translation[13] = 111_01101000000000000000000
w[13] = 2 * (w[12] - q[13] * D) = 2 * (
	111_00000010000000000000000 +
	001_01010110000000000000000
) = 2 * 000_01011000000000000000000 = 
000_10110000000000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 001111111111111110000011 = 4194179
D[WIDTH-1:0] = 000000000010000000110000 = 8240
Q[WIDTH-1:0] = X / D = 509 = 000000000000000111111101
REM[WIDTH-1:0] = 4194179 - 8240 * 509 = 19 = 000000000000000000010011

CLZ_X = 2
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 8
迭代次数:
iter_num = CLZ_DIFF + 1 = 9
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111111111111111000001100
Divisor[WIDTH-1:0] 		= 100000001100000000000000

+ D[(WIDTH + 2)-1:0] = 001_00000001100000000000000
+2D[(WIDTH + 2)-1:0] = 010_00000011000000000000000
- D[(WIDTH + 2)-1:0] = 110_11111110100000000000000
-2D[(WIDTH + 2)-1:0] = 101_11111101000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[9] = 010_00000100001100000000000 >= 0;
(w[final] / 2) + (-D) = 001_00000010000110000000000 + 110_11111110100000000000000 = 
00000000000100110000000000 >= 0 -> (w[final] / 2) "belongs to [+D, +2D)";
// 最后一次迭代的商
q_pos = 1111_1110_0
q_neg = 0000_0000_0

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 111111100;
(w[final] / 2) "belongs to [+D, +2D)" -> quotient_correction_coefficient = 1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 111111101;

(w[final] / 2) "belongs to [+D, +2D)" -> remainder_correction_coefficient = 1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
(001_00000010000110000000000 + 110_11111110100000000000000) >> 10 = 
000000000100110000000000 >> 10
000000000000000000010011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 001111111111111110000011 = 4194179
D[WIDTH-1:0] = 000000001000000011000000 = 32960
Q[WIDTH-1:0] = X / D = 127 = 000000000000000001111111
REM[WIDTH-1:0] = 4194179 - 32960 * 127 = 8259 = 000000000010000001000011

CLZ_X = 2
CLZ_D = 8
CLZ_DIFF = CLZ_D - CLZ_X = 6
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 8
q[7] = +2
q[8] = +1
q_pos = 1111_1101
q_neg = 0000_0000
q_pos - q_neg = 11111101
w[8] = 011_00000101000110000000000 >= 0
w[8] / 2 = 001_10000010100011000000000
001_10000010100011000000000 + (-D) = 
001_10000010100011000000000 + 110_11111110100000000000000 = 
000_10000001000011000000000

010000001000011000000000 >> (CLZ_D + 1) = 
000000000010000001000011

// ---------------------------------------------------------------------------------------------------------------------------------------







初始化:
w[0][(WIDTH + 2)-1:0] =  001_11111111111111000001100
w_sum_translation[0] = w_sum[0] =  001_11111111111111000001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_11111111111110000011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11111101000000000000000
w_sum_translation[1] = 001_11111111111110000011000
w_carry_translation[1] = 111_11111101000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11111111111111000001100 +
	110_11111110100000000000000
) = 2 * 000_11111110011111000001100 = 
001_11111100111110000011000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_11111111111100000110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11111010000000000000000
w_sum_translation[2] = 001_11111111111100000110000
w_carry_translation[2] = 001_11111010000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_01 -> q[3] = +2
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	001_11111100111110000011000 +
	000_00000000000000000000000
) = 2 * 001_11111100111110000011000 = 
011_11111001111100000110000
q_pos = 110
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_11110001111000001100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11111100000000000000000
w_sum_translation[3] = 001_11110001111000001100000
w_carry_translation[3] = 001_11111100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_01 -> q[4] = +2
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	011_11111001111100000110000 +
	101_11111101000000000000000
) = 2 * 001_11110110111100000110000 = 
011_11101101111000001100000
q_pos = 1110
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_11100001110000011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11110100000000000000000
w_sum_translation[4] = 001_11100001110000011000000
w_carry_translation[4] = 001_11110100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[5] = +2
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	011_11101101111000001100000 +
	101_11111101000000000000000
) = 2 * 001_11101010111000001100000 = 
011_11010101110000011000000
q_pos = 1111_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_11010001100000110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11010100000000000000000
w_sum_translation[5] = 001_11010001100000110000000
w_carry_translation[5] = 001_11010100000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	011_11010101110000011000000 +
	101_11111101000000000000000
) = 2 * 001_11010010110000011000000 = 
011_10100101100000110000000
q_pos = 1111_10
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_11110001000001100000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_01010100000000000000000
w_sum_translation[6] = 001_11110001000001100000000
w_carry_translation[6] = 001_01010100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_01 -> q[7] = +2
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_10100101100000110000000 +
	101_11111101000000000000000
) = 2 * 001_10100010100000110000000 = 
011_01000101000001100000000
q_pos = 1111_110
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_10110000000011000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_11010100000000000000000
w_sum_translation[7] = 000_10110000000011000000000
w_carry_translation[7] = 001_11010100000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	011_01000101000001100000000 +
	101_11111101000000000000000
) = 2 * 001_01000010000001100000000 = 
010_10000100000011000000000
q_pos = 1111_1101
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
111_00110101000110000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
011_11010000000000000000000
w_sum_translation[8] = 001_00110101000110000000000
w_carry_translation[8] = 001_11010000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 01_01 -> q[9] = +2
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_10000100000011000000000 +
	110_11111110100000000000000
) = 2 * 001_10000010100011000000000 = 
011_00000101000110000000000
q_pos = 1111_1110_0
q_neg = 0000_0000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_00110000001100000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
011_11010100000000000000000
w_sum_translation[9] = 000_00110000001100000000000
w_carry_translation[9] = 001_11010100000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_01 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	011_00000101000110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000010000110000000000 = 
010_00000100001100000000000
q_pos = 1111_1110_01
q_neg = 0000_0000_00



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 001000000010011111110011 = 2107379
D[WIDTH-1:0] = 001111111100001100000000 = 4178688
Q[WIDTH-1:0] = X / D = 0 = 000000000000000000000000
REM[WIDTH-1:0] = 2107379 - 4178688 * 0 = 2107379 = 001000000010011111110011

CLZ_X = 2
CLZ_D = 2
CLZ_DIFF = CLZ_D - CLZ_X = 0
迭代次数:
iter_num = CLZ_DIFF + 1 = 1
规格化操作之后:
Dividend[WIDTH-1:0] 	= 100000001001111111001100
Divisor[WIDTH-1:0] 		= 111111110000110000000000

+ D[(WIDTH + 2)-1:0] = 001_11111110000110000000000
+2D[(WIDTH + 2)-1:0] = 011_11111100001100000000000
- D[(WIDTH + 2)-1:0] = 110_00000001111010000000000
-2D[(WIDTH + 2)-1:0] = 100_00000011110100000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[1] = 110_00000110010011110011000 < 0;
(w[final] / 2) + (D) = 111_00000011001001111001100 + 001_11111110000110000000000 = 
00100000001001111111001100 >= 0 -> (w[final] / 2) "belongs to [-D, +0)";
// 最后一次迭代的商
q_pos = 1
q_neg = 0

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 1;
(w[final] / 2) "belongs to [-D, +0)" -> quotient_correction_coefficient = -1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 0;

(w[final] / 2) "belongs to [-D, +0)" -> remainder_correction_coefficient = -1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
(111_00000011001001111001100 + 001_11111110000110000000000) >> 2 = 
100000001001111111001100 >> 2
001000000010011111110011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 余数是负数
REM[WIDTH-1:0] = -2107379 = 110111111101100000001101

w_sum_translation[final] = 000_00000010011111110011000
w_carry_translation[final] = 110_00000011110100000000000
~w_sum_translation[final] = 111_11111101100000001100111
~w_carry_translation[final] = 001_11111100001011111111111

w[final] = ~w_sum_translation[final] + ~w_carry_translation[final] + 2'b10 = 001_11111001101100001101000 >= 0
(w[final] / 2) + (-D) = 000_11111100110110000110100 + 110_00000001111010000000000 = 
110_11111110110000000110100 < 0 -> (w[final] / 2) "belongs to (0, +D]".

remainder_calculated[WIDTH-1:0] = ((w[final] / 2) + (-D)) >> CLZ_D = 
(000_11111100110110000110100 + 110_00000001111010000000000) >> 2 = 
110_11111110110000000110100 >> 2 = 
110111111101100000001101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_00000001001111111001100
w_sum_translation[0] = w_sum[0] =  001_00000001001111111001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_00000010011111110011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_00000011110100000000000
w_sum_translation[1] = 000_00000010011111110011000
w_carry_translation[1] = 110_00000011110100000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_00000001001111111001100 +
	110_00000001111010000000000
) = 2 * 111_00000011001001111001100 = 
110_00000110010011110011000
q_pos = 10
q_neg = 00


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000000111101001111111000 = 250872
D[WIDTH-1:0] = 000000000000000010111010 = 186
Q[WIDTH-1:0] = X / D = 1348 = 000000000000010101000100
REM[WIDTH-1:0] = 250872 - 186 * 1348 = 144 = 000000000000000010010000

CLZ_X = 6
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 10
迭代次数:
iter_num = CLZ_DIFF + 1 = 11
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111101001111111000000000
Divisor[WIDTH-1:0] 		= 101110100000000000000000

+ D[(WIDTH + 2)-1:0] = 001_01110100000000000000000
+2D[(WIDTH + 2)-1:0] = 010_11101000000000000000000
- D[(WIDTH + 2)-1:0] = 110_10001100000000000000000
-2D[(WIDTH + 2)-1:0] = 101_00011000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[11] = 111_01011000000000000000000 < 0;
(w[final] / 2) + (D) = 111_10101100000000000000000 + 001_01110100000000000000000 = 
00100100000000000000000000 >= 0 -> (w[final] / 2) "belongs to [-D, +0)";
// 最后一次迭代的商
q_pos = 1011_0000_110
q_neg = 0000_1000_001

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 010101000101;
(w[final] / 2) "belongs to [-D, +0)" -> quotient_correction_coefficient = -1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 010101000100;

(w[final] / 2) "belongs to [-D, +0)" -> remainder_correction_coefficient = -1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
(111_10101100000000000000000 + 001_01110100000000000000000) >> 16 = 
100100000000000000000000 >> 16
000000000000000010010000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_11101001111111000000000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_11010011111110000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_00011000000000000000000
w_sum_translation[1] = 001_11010011111110000000000
w_carry_translation[1] = 111_00011000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11101001111111000000000 +
	110_10001100000000000000000
) = 2 * 000_01110101111111000000000 = 
000_11101011111110000000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_10100111111100000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_00110000000000000000000
w_sum_translation[2] = 001_10100111111100000000000
w_carry_translation[2] = 000_00110000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_00 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_11101011111110000000000 +
	000_00000000000000000000000
) = 2 * 000_11101011111110000000000 = 
001_11010111111100000000000
q_pos = 101
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_00110111111000000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_10010000000000000000000
w_sum_translation[3] = 000_00110111111000000000000
w_carry_translation[3] = 000_10010000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_00 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_11010111111100000000000 +
	110_10001100000000000000000
) = 2 * 000_01100011111100000000000 = 
000_11000111111000000000000
q_pos = 1011
q_neg = 0000


w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_01010111110000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_01010000000000000000000
w_sum_translation[4] = 000_01010111110000000000000
w_carry_translation[4] = 110_01010000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_11000111111000000000000 +
	110_10001100000000000000000
) = 2 * 111_01010011111000000000000 = 
110_10100111110000000000000
q_pos = 1011_0
q_neg = 0000_0
abs(w[4]) = 001_01011000010000000000000
+D = 001_01110100000000000000000

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_10101111100000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_10100000000000000000000
w_sum_translation[5] = 110_10101111100000000000000
w_carry_translation[5] = 110_10100000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 10_10 -> q[6] = -2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	110_10100111110000000000000 +
	000_00000000000000000000000
) = 2 * 110_10100111110000000000000 = 
101_01001111100000000000000
q_pos = 1011_00
q_neg = 0000_10

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_11001111000000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_10100000000000000000000
w_sum_translation[6] = 111_11001111000000000000000
w_carry_translation[6] = 000_10100000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 11_00 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	101_01001111100000000000000 +
	010_11101000000000000000000
) = 2 * 000_00110111100000000000000 = 
000_01101111000000000000000
q_pos = 1011_000
q_neg = 0000_100

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_10011110000000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
001_01000000000000000000000
w_sum_translation[7] = 111_10011110000000000000000
w_carry_translation[7] = 001_01000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 11_01 -> q[8] = 0
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_01101111000000000000000 +
	000_00000000000000000000000
) = 2 * 000_01101111000000000000000 = 
000_11011110000000000000000
q_pos = 1011_0000
q_neg = 0000_1000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
111_00111100000000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
010_10000000000000000000000
w_sum_translation[8] = 001_00111100000000000000000
w_carry_translation[8] = 000_10000000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 01_00 -> q[9] = +1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	000_11011110000000000000000 +
	000_00000000000000000000000
) = 2 * 000_11011110000000000000000 = 
001_10111100000000000000000
q_pos = 1011_0000_1
q_neg = 0000_1000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
010_01100000000000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_00110000000000000000000
w_sum_translation[9] = 000_01100000000000000000000
w_carry_translation[9] = 000_00110000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_00 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	001_10111100000000000000000 +
	110_10001100000000000000000
) = 2 * 000_01001000000000000000000 = 
000_10010000000000000000000
q_pos = 1011_0000_11
q_neg = 0000_1000_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_10111000000000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
100_10000000000000000000000
w_sum_translation[10] = 111_10111000000000000000000
w_carry_translation[10] = 110_10000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 11_10 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	000_10010000000000000000000 +
	110_10001100000000000000000
) = 2 * 111_00011100000000000000000 = 
110_00111000000000000000000
q_pos = 1011_0000_110
q_neg = 0000_1000_001

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_10011000000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
010_11000000000000000000000
w_sum_translation[11] = 110_10011000000000000000000
w_carry_translation[11] = 000_11000000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_00 -> q[12] = 0
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	110_00111000000000000000000 +
	001_01110100000000000000000
) = 2 * 111_10101100000000000000000 = 
111_01011000000000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000111011110000111101110 = 1958382
D[WIDTH-1:0] = 000000000011101101000000 = 15168
Q[WIDTH-1:0] = X / D = 129 = 000000000000000010000001
REM[WIDTH-1:0] = 1958382 - 15168 * 129 = 1710 = 000000000000011010101110

CLZ_X = 3
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 7
迭代次数
iter_num = CLZ_DIFF + 1 = 8
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111011110000111101110000
Divisor[WIDTH-1:0] 		= 111011010000000000000000

+ D[(WIDTH + 2)-1:0] = 001_11011010000000000000000
+2D[(WIDTH + 2)-1:0] = 011_10110100000000000000000
- D[(WIDTH + 2)-1:0] = 110_00100110000000000000000
-2D[(WIDTH + 2)-1:0] = 100_01001100000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8] = 100_10110110111000000000000 < 0;
(w[final] / 2) + (D) = 110_01011011011100000000000 + 001_11011010000000000000000 = 
00000110101011100000000000 >= 0 -> (w[final] / 2) "belongs to [-D, +0)";
// 最后一次迭代的商
q_pos = 1000_0010
q_neg = 0000_0000

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 10000010;
(w[final] / 2) "belongs to [-D, +0)" -> quotient_correction_coefficient = -1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 10000001;

(w[final] / 2) "belongs to [-D, +0)" -> remainder_correction_coefficient = -1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
(110_01011011011100000000000 + 001_11011010000000000000000) >> 10 = 
000110101011100000000000 >> 10
000000000000011010101110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_11011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_11011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_10111100001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_01001100000000000000000
w_sum_translation[1] = 001_10111100001111011100000
w_carry_translation[1] = 110_01001100000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11011110000111101110000 +
	110_00100110000000000000000
) = 2 * 000_00000100000111101110000 = 
000_00001000001111011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_01111000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_10011000000000000000000
w_sum_translation[2] = 001_01111000011110111000000
w_carry_translation[2] = 110_10011000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_00001000001111011100000 +
	000_00000000000000000000000
) = 2 * 000_00001000001111011100000 = 
000_00010000011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_11110000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
101_00110000000000000000000
w_sum_translation[3] = 000_11110000111101110000000
w_carry_translation[3] = 111_00110000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00010000011110111000000 +
	000_00000000000000000000000
) = 2 * 000_00010000011110111000000 = 
000_00100000111101110000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_11100001111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_01100000000000000000000
w_sum_translation[4] = 001_11100001111011100000000
w_carry_translation[4] = 110_01100000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00100000111101110000000 +
	000_00000000000000000000000
) = 2 * 000_00100000111101110000000 = 
000_01000001111011100000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11000011110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_11000000000000000000000
w_sum_translation[5] = 001_11000011110111000000000
w_carry_translation[5] = 110_11000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_01000001111011100000000 +
	000_00000000000000000000000
) = 2 * 000_01000001111011100000000 = 
000_10000011110111000000000
q_pos = 1000_00
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_10000111101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_10000000000000000000000
w_sum_translation[6] = 001_10000111101110000000000
w_carry_translation[6] = 111_10000000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_11 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_10000011110111000000000 +
	000_00000000000000000000000
) = 2 * 000_10000011110111000000000 = 
001_00000111101110000000000
q_pos = 1000_000
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_00001111011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_00000000000000000000000
w_sum_translation[7] = 001_00001111011100000000000
w_carry_translation[7] = 001_00000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 01_01 -> q[8] = +2
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	001_00000111101110000000000 +
	000_00000000000000000000000
) = 2 * 001_00000111101110000000000 = 
010_00001111011100000000000
q_pos = 1000_0010
q_neg = 0000_0000

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_00001111011100000000000 +
	100_01001100000000000000000
) = 2 * 110_01011011011100000000000 = 
100_10110110111000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000010001100010111011110011 = 4599539
D[WIDTH-1:0] = 0000000000000001000111010100 = 4564
Q[WIDTH-1:0] = X / D = 1007 = 0000000000000000001111101111
REM[WIDTH-1:0] = 4599539 - 4564 * 1007 = 3591 = 0000000000000000111000000111

CLZ_X = 5
CLZ_D = 15
CLZ_DIFF = CLZ_D - CLZ_X = 10
迭代次数:
iter_num = CLZ_DIFF + 1 = 11
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000110001011101111001100000
Divisor[WIDTH-1:0] 		= 1000111010100000000000000000

+ D[(WIDTH + 2)-1:0] = 001_000111010100000000000000000
+2D[(WIDTH + 2)-1:0] = 010_001110101000000000000000000
- D[(WIDTH + 2)-1:0] = 110_111000101100000000000000000
-2D[(WIDTH + 2)-1:0] = 101_110001011000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[11] = 101_010010111110000000000000000 < 0;
(w[final] / 2) + (D) = 110_101001011111000000000000000 + 001_000111010100000000000000000 = 
111110000110011000000000000000 < 0 -> (w[final] / 2) "belongs to [-2D, -D)";
// 最后一次迭代的商
q_pos = 1000_0000_000
q_neg = 0000_0001_111

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 001111110001;
(w[final] / 2) "belongs to [-2D, -D)" -> quotient_correction_coefficient = -2;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 001111101111;

(w[final] / 2) "belongs to [-2D, -D)" -> remainder_correction_coefficient = -2;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[0 +: WIDTH]) >> CLZ_D = 
(110_101001011111000000000000000 + 010_001110101000000000000000000) >> 15 = 
0111000000111000000000000000 >> 15
0000000000000000111000000111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 余数是负数
REM[WIDTH-1:0] = -3591 = 1111111111111111000111111001

w_sum_translation[final] = 110_111110111110000000000000000
w_carry_translation[final] = 110_010100000000000000000000000
~w_sum_translation[final] = 001_000001000001111111111111111
~w_carry_translation[final] = 001_101011111111111111111111111

w[final] = ~w_sum_translation[final] + ~w_carry_translation[final] + 2'b10 = 010_101101000010000000000000000 >= 0
(w[final] / 2) + (-D) = 001_010110100001000000000000000 + 110_111000101100000000000000000 = 
000_001111001101000000000000000 >= 0 -> (w[final] / 2) "belongs to (+D, +2D]".

remainder_calculated[WIDTH-1:0] = ((w[final] / 2) + -2D) >> CLZ_D = 
(001_010110100001000000000000000 + 101_110001011000000000000000000) >> 15 = 
111_000111111001000000000000000 >> 15 = 
1111111111111111000111111001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 0000010001100010111011110011 = 4599539
D[WIDTH-1:0] = 0000000000010001110101000000 = 73024
Q[WIDTH-1:0] = X / D = 62 = 0000000000000000000000111110
REM[WIDTH-1:0] = 4599539 - 73024 * 62 = 72051 = 0000000000010001100101110011

CLZ_X = 5
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 6
迭代次数:
iter_num = CLZ_DIFF + 2 = 8
q[8] = -1
q_pos = 1000_0000
q_neg = 0000_0001
q_pos - q_neg = 01111111

w[8] = 101_101101100100110000000000000 < 0
w[8] / 2 = 110_110110110010011000000000000
110_110110110010011000000000000 + (D) = 
110_110110110010011000000000000 + 001_000111010100000000000000000 = 
111_111110000110011000000000000

111_111110000110011000000000000 + (D) = 
001_000101011010011000000000000

1000101011010011000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------



初始化:
w[0][(WIDTH + 2)-1:0] =  001_000110001011101111001100000
w_sum_translation[0] = w_sum[0] =  001_000110001011101111001100000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_001100010111011110011000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_110001011000000000000000000
w_sum_translation[1] = 000_001100010111011110011000000
w_carry_translation[1] = 111_110001011000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_000110001011101111001100000 +
	110_111000101100000000000000000
) = 2 * 111_111110110111101111001100000 = 
111_111101101111011110011000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_011000101110111100110000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_100010110000000000000000000
w_sum_translation[2] = 000_011000101110111100110000000
w_carry_translation[2] = 111_100010110000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	111_111101101111011110011000000 +
	000_000000000000000000000000000
) = 2 * 111_111101101111011110011000000 = 
111_111011011110111100110000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_110001011101111001100000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_000101100000000000000000000
w_sum_translation[3] = 000_110001011101111001100000000
w_carry_translation[3] = 111_000101100000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	111_111011011110111100110000000 +
	000_000000000000000000000000000
) = 2 * 111_111011011110111100110000000 = 
111_110110111101111001100000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_100010111011110011000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_001011000000000000000000000
w_sum_translation[4] = 001_100010111011110011000000000
w_carry_translation[4] = 110_001011000000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	111_110110111101111001100000000 +
	000_000000000000000000000000000
) = 2 * 111_110110111101111001100000000 = 
111_101101111011110011000000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_000101110111100110000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_010110000000000000000000000
w_sum_translation[5] = 001_000101110111100110000000000
w_carry_translation[5] = 110_010110000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	111_101101111011110011000000000 +
	000_000000000000000000000000000
) = 2 * 111_101101111011110011000000000 = 
111_011011110111100110000000000
q_pos = 1000_00
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_001011101111001100000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
100_101100000000000000000000000
w_sum_translation[6] = 000_001011101111001100000000000
w_carry_translation[6] = 110_101100000000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 00_10 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	111_011011110111100110000000000 +
	000_000000000000000000000000000
) = 2 * 111_011011110111100110000000000 = 
110_110111101111001100000000000
q_pos = 1000_000
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
000_010111011110011000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
101_011000000000000000000000000
w_sum_translation[7] = 110_010111011110011000000000000
w_carry_translation[7] = 111_011000000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 10_11 -> q[8] = -1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	110_110111101111001100000000000 +
	000_000000000000000000000000000
) = 2 * 110_110111101111001100000000000 = 
101_101111011110011000000000000
q_pos = 1000_0000
q_neg = 0000_0001


w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
000_010000010100110000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
101_011101010000000000000000000
w_sum_translation[8] = 110_010000010100110000000000000
w_carry_translation[8] = 111_011101010000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_11 -> q[9] = -1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	101_101111011110011000000000000 +
	001_000111010100000000000000000
) = 2 * 110_110110110010011000000000000 = 
101_101101100100110000000000000
q_pos = 1000_0000_0
q_neg = 0000_0001_1

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
000_010100100001100000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
101_010101010000000000000000000
w_sum_translation[9] = 110_010100100001100000000000000
w_carry_translation[9] = 111_010101010000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_11 -> q[10] = -1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	101_101101100100110000000000000 +
	001_000111010100000000000000000
) = 2 * 110_110100111000110000000000000 = 
101_101001110001100000000000000
q_pos = 1000_0000_00
q_neg = 0000_0001_11

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
000_001101001011000000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
101_010101000000000000000000000
w_sum_translation[10] = 110_001101001011000000000000000
w_carry_translation[10] = 111_010101000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 10_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	101_101001110001100000000000000 +
	001_000111010100000000000000000
) = 2 * 110_110001000101100000000000000 = 
101_100010001011000000000000000
q_pos = 1000_0000_000
q_neg = 0000_0001_111

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
000_111110111110000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_010100000000000000000000000
w_sum_translation[11] = 110_111110111110000000000000000
w_carry_translation[11] = 110_010100000000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_10 -> q[12] = -2
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	101_100010001011000000000000000 +
	001_000111010100000000000000000
) = 2 * 110_101001011111000000000000000 = 
101_010010111110000000000000000



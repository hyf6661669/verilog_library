



a = 0.10010001111
b = 0.10000010001
a / b = 1.00011110111111000100111110101101010111110010101110
a_scaled = a << 1 = 1.00100011110000
b_scaled = b << 1 = 1.00000100010000

d   = 00100000100010000
2d  = 01000001000100000
~d  = 11011111011101111
~2d = 10111110111011111
-d  = 11011111011110000
-2d = 10111110111100000

// ==================================================================================================
rem_init = 00001001000111100
rem_s[0] = rem_init = 00001001000111100
rem_c[0] = 00000000000000000
rem[0] = 00001001000111100

// ================
// BigIter[0]
d   = 00100000100010000
2d  = 01000001000100000
~d  = 11011111011101111
~2d = 10111110111011111
-d  = 11011111011110000
-2d = 10111110111100000
// ================
// stage[0]
rem_s[0][14:9] + rem_c[0][14:9] = 
001001 + 
000000 = 
001001, belongs to "[4/8, 12/8]" -> q[0] = +1
q_pos = 01
q_neg = 00
q_pos - q_neg = 01
a / b = 1.00011110111111000100111110101101010111110010101110

// stage[1]
rem_s[1] = 00100100011110000
rem_c[1] = 11011111011110000
-> 
rem[1] = 
00100100011110000 + 
11011111011110000 = 
00000011111100000

rem_s[1][14:9] + rem_c[1][14:9] = 
100100 + 
011111 = 
000011, belongs to "[-3/8, 3/8]" -> q[1] = 0
q_pos = 0100
q_neg = 0000
q_pos - q_neg = 0100
a / b = 1.00011110111111000100111110101101010111110010101110

// TODO
adder_9b = (rem_s[1] << 2)[16:8] + (rem_c[1] << 2)[16:8] = 
100100011 + 
011111011 =
000011110
adder_9b[8:3] = 000011, 此时adder_9b[3].carry = 0, 按照TABLE II(b), 应该选择q[1] = +1
->
q_pos = 0101
q_neg = 0000
q_pos - q_neg = 0101
a / b = 1.00011110111111000100111110101101010111110010101110
1.000110

// stage[2]
rem_s[2] = 11110111010011000
rem_c[2] = 00000001011001000
->
rem[2] = 
10110000110000000 + 
01000111111100000 = 
11111000101100000

rem_s[2][14:9] + rem_c[2][14:9] = 
110111 + 
000001 = 
111000, belongs to "[-12/8, -5/8]" -> q[2] = -1
q_pos = 100000
q_neg = 001001
q_pos - q_neg = 010111
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[1] * d) << 2)[16:10] + adder_9b[6:0]
0001111 +
1100001 = 
1110000, adder_7b[6:1] = 111000, belongs to "[-12/8, -4/8]" -> q[2] = -1
测试"WIDTH = 16"时, 使用"WIDTH = 32"的计算模块进行SRT迭代的设计.

// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 16;
ITN = InTerNal
ITN_W = 1 + (2 * WIDTH) = 33;
0_00000000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0001010010010100 = 5268
D[WIDTH-1:0] = 0000001000000011 = 515
Q[WIDTH-1:0] = X / D = 10 = 0000000000001010
REM[WIDTH-1:0] = 5268 - 515 * 10 = 118 = 0000000001110110

CLZ_X = 3
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 3
Normalized_D = 1000000011000000
根据D的值, 可得选择常数:
m[-1] = -13
m[ 0] = - 4
m[+1] = + 4
m[+2] = +12

+ D[ITN_W-1:0] = 0_10000000110000000000000000000000
+2D[ITN_W-1:0] = 1_00000001100000000000000000000000
- D[ITN_W-1:0] = 1_01111111010000000000000000000000
-2D[ITN_W-1:0] = 0_11111110100000000000000000000000

l_shift_num = CLZ_D = 6
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000000001010010010100 << 6 = 
0_00000000000001010010010100000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:0] = 0_00000000000001010010010100000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w[1] = w[0] << 2 - q[1] * D = 
0_00000000000101001001010000000000 + 
0_00000000000000000000000000000000 = 
0_00000000000101001001010000000000
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
w[2] = w[1] << 2 - q[2] * D = 
0_00000000010100100101000000000000 + 
0_00000000000000000000000000000000 = 
0_00000000010100100101000000000000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00

ITER[2]:
w[3] = w[2] << 2 - q[3] * D = 
0_00000001010010010100000000000000 + 
0_00000000000000000000000000000000 = 
0_00000001010010010100000000000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000

ITER[3]:
w[4] = w[3] << 2 - q[4] * D = 
0_00000101001001010000000000000000 + 
0_00000000000000000000000000000000 = 
0_00000101001001010000000000000000
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00

ITER[4]:
w[5] = w[4] << 2 - q[5] * D = 
0_00010100100101000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00010100100101000000000000000000
(4 * w[5])_trunc_3_4 = 000_0101, "belongs to [m[+1], m[+2])" -> q[6] = +1
q_pos = 0000_0000_0001
q_neg = 0000_0000_0000

ITER[5]:
w[6] = w[5] << 2 - q[6] * D = 
0_01010010010100000000000000000000 + 
1_01111111010000000000000000000000 = 
1_11010001100100000000000000000000
(4 * w[6])_trunc_3_4 = 111_0100, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0000_0000_0001_00
q_neg = 0000_0000_0000_01

ITER[6]:
w[7] = w[6] << 2 - q[7] * D = 
1_01000110010000000000000000000000 + 
0_10000000110000000000000000000000 = 
1_11000111000000000000000000000000
(4 * w[7])_trunc_3_4 = 111_0001, "belongs to [-Inf, m[-1])" -> q[8] = -2
q_pos = 0000_0000_0001_0000
q_neg = 0000_0000_0000_0110

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[8] = w[7] << 2 - q[8] * D = 
1_00011100000000000000000000000000 + 
1_00000001100000000000000000000000 = 
0_00011101100000000000000000000000 >= 0

rem = (w[8])_reduced >> CLZ_D = 
0001110110000000 >> 6
0000000001110110

q_final = corr(q_pos - q_neg) = 0000000000001010
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110011110101 = 3317
D[WIDTH-1:0] = 0000000000000011 = 3
Q[WIDTH-1:0] = X / D = 1105 = 0000010001010001
REM[WIDTH-1:0] = 3317 - 3 * 1105 = 2 = 0000000000000010

CLZ_X = 4
CLZ_D = 14
CLZ_DIFF = CLZ_D - CLZ_X = 10
Normalized_D = 1100000000000000
根据D的值, 可得选择常数:
m[-1] = -18
m[ 0] = - 6
m[+1] = + 6
m[+2] = +18

+ D[ITN_W-1:0] = 0_11000000000000000000000000000000
+2D[ITN_W-1:0] = 1_10000000000000000000000000000000
- D[ITN_W-1:0] = 1_01000000000000000000000000000000
-2D[ITN_W-1:0] = 0_10000000000000000000000000000000

l_shift_num = CLZ_D = 14
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000000000110011110101 << 14 = 
0_00000011001111010100000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:0] = 0_00000011001111010100000000000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w[1] = w[0] << 2 - q[1] * D = 
0_00001100111101010000000000000000 + 
0_00000000000000000000000000000000 = 
0_00001100111101010000000000000000
(4 * w[1])_trunc_3_4 = 000_0011, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
w[2] = w[1] << 2 - q[2] * D = 
0_00110011110101000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00110011110101000000000000000000
(4 * w[2])_trunc_3_4 = 000_1100, "belongs to [m[+1], m[+2])" -> q[3] = +1
q_pos = 0000_01
q_neg = 0000_00

ITER[2]:
w[3] = w[2] << 2 - q[3] * D = 
0_11001111010100000000000000000000 + 
1_01000000000000000000000000000000 = 
0_00001111010100000000000000000000
(4 * w[3])_trunc_3_4 = 000_0011, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0100
q_neg = 0000_0000

ITER[3]:
w[4] = w[3] << 2 - q[4] * D = 
0_00111101010000000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00111101010000000000000000000000
(4 * w[4])_trunc_3_4 = 000_1111, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0000_0100_01
q_neg = 0000_0000_00

ITER[4]:
w[5] = w[4] << 2 - q[5] * D = 
0_11110101000000000000000000000000 + 
1_01000000000000000000000000000000 = 
0_00110101000000000000000000000000
(4 * w[5])_trunc_3_4 = 000_1101, "belongs to [m[+1], m[+2])" -> q[6] = +1
q_pos = 0000_0100_0101
q_neg = 0000_0000_0000

ITER[5]:
w[6] = w[5] << 2 - q[6] * D = 
0_11010100000000000000000000000000 + 
1_01000000000000000000000000000000 = 
0_00010100000000000000000000000000
(4 * w[6])_trunc_3_4 = 000_0101, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0100_0101_00
q_neg = 0000_0000_0000_00

ITER[6]:
w[7] = w[6] << 2 - q[7] * D = 
0_01010000000000000000000000000000 + 
0_00000000000000000000000000000000 = 
0_01010000000000000000000000000000
(4 * w[7])_trunc_3_4 = 001_0100, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0000_0100_0101_0010
q_neg = 0000_0000_0000_0000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[8] = w[7] << 2 - q[8] * D = 
1_01000000000000000000000000000000 + 
0_10000000000000000000000000000000 = 
1_11000000000000000000000000000000 < 0

rem = (w[8] + D)_reduced >> CLZ_D = 
(11000000000000000000000000000000 + 11000000000000000000000000000000)_reduced >> 14
1000000000000000 >> 14 = 
0000000000000010

q_final = corr(q_pos - q_neg) = 0000010001010001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000000010011101 = 157
D[WIDTH-1:0] = 0000111000010010 = 3602
Q[WIDTH-1:0] = X / D = 0 = 0000000000000000
REM[WIDTH-1:0] = 157 - 3602 * 0 = 157 = 0000000010011101

CLZ_X = 8
CLZ_D = 4
CLZ_DIFF = CLZ_D - CLZ_X = -4
Normalized_D = 1110000100100000
根据D的值, 可得选择常数:
m[-1] = -22
m[ 0] = - 8
m[+1] = + 8
m[+2] = +22

+ D[ITN_W-1:0] = 0_11100001001000000000000000000000
+2D[ITN_W-1:0] = 1_11000010010000000000000000000000
- D[ITN_W-1:0] = 1_00011110111000000000000000000000
-2D[ITN_W-1:0] = 0_00111101110000000000000000000000

l_shift_num = CLZ_D = 4
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000000000000010011101 << 4 = 
0_00000000000000000000100111010000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:0] = 0_00000000000000000000100111010000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w[1] = w[0] << 2 - q[1] * D = 
0_00000000000000000010011101000000 + 
0_00000000000000000000000000000000 = 
0_00000000000000000010011101000000
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
w[2] = w[1] << 2 - q[2] * D = 
0_00000000000000001001110100000000 + 
0_00000000000000000000000000000000 = 
0_00000000000000001001110100000000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00

ITER[2]:
w[3] = w[2] << 2 - q[3] * D = 
0_00000000000000100111010000000000 + 
0_00000000000000000000000000000000 = 
0_00000000000000100111010000000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000

ITER[3]:
w[4] = w[3] << 2 - q[4] * D = 
0_00000000000010011101000000000000 + 
0_00000000000000000000000000000000 = 
0_00000000000010011101000000000000
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00

ITER[4]:
w[5] = w[4] << 2 - q[5] * D = 
0_00000000001001110100000000000000 + 
0_00000000000000000000000000000000 = 
0_00000000001001110100000000000000
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000

ITER[5]:
w[6] = w[5] << 2 - q[6] * D = 
0_00000000100111010000000000000000 + 
0_00000000000000000000000000000000 = 
0_00000000100111010000000000000000
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00

ITER[6]:
w[7] = w[6] << 2 - q[7] * D = 
0_00000010011101000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00000010011101000000000000000000
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[8] = w[7] << 2 - q[8] * D = 
0_00001001110100000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00001001110100000000000000000000 >= 0

rem = (w[8])_reduced >> CLZ_D = 
0000100111010000 >> 4 = 
0000000010011101

q_final = corr(q_pos - q_neg) = 0000000000000000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------



// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 16;
ITN = InTerNal
ITN_W = 1 + WIDTH = 17;
0_0000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1010100110100011
D[WIDTH-1:0] = 0110101101111101
Q[WIDTH-1:0] = X / D = 0000000000000000
REM[WIDTH-1:0] = 0011111000100110

CLZ_X = 0
CLZ_D = 1
CLZ_DIFF = CLZ_D - CLZ_X = 1
Normalized_D = 1101011011111010
根据D的值, 可得选择常数:
m[-1] = -20
m[ 0] = - 8
m[+1] = + 6
m[+2] = +20

+ D[ITN_W-1:0] = 0_1101011011111010
+2D[ITN_W-1:0] = 1_1010110111110100
- D[ITN_W-1:0] = 1_0010100100000110
-2D[ITN_W-1:0] = 0_0101001000001100
~2D[ITN_W-1:0] = 0_0101001000001011

l_shift_num = CLZ_D = 1
shifted_dividend[(2 * WIDTH + 1)-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000001010100110100011 << 1 = 
0_00000000000000010101001101000110

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:0] = 0_0000000000000001
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
0101001101000110

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_0000000000000101 + 
0_0000000000000000 = 
0_0000000000000101
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1][WIDTH-1:0] = temp_dividend[0][WIDTH-1:0] << 2 = 
0100110100011000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_0000000000010101 + 
0_0000000000000000 = 
0_0000000000010101
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2][WIDTH-1:0] = temp_dividend[1][WIDTH-1:0] << 2 = 
0011010001100000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_0000000001010100 + 
0_0000000000000000 = 
0_0000000001010100
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3][WIDTH-1:0] = temp_dividend[2][WIDTH-1:0] << 2 = 
1101000110000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_0000000101010011 + 
0_0000000000000000 = 
0_0000000101010011
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4][WIDTH-1:0] = temp_dividend[3][WIDTH-1:0] << 2 = 
0100011000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_0000010101001101 + 
0_0000000000000000 = 
0_0000010101001101
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5][WIDTH-1:0] = temp_dividend[4][WIDTH-1:0] << 2 = 
0001100000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_0001010100110100 + 
0_0000000000000000 = 
0_0001010100110100
(4 * w[6])_trunc_3_4 = 000_0101, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6][WIDTH-1:0] = temp_dividend[5][WIDTH-1:0] << 2 = 
0110000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_0101010011010001 + 
0_0000000000000000 = 
0_0101010011010001
(4 * w[7])_trunc_3_4 = 001_0101, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0000_0000_0000_0010
q_neg = 0000_0000_0000_0000
temp_dividend[7][WIDTH-1:0] = temp_dividend[6][WIDTH-1:0] << 2 = 
1000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
1_0101001101000110 + 
0_0101001000001100 = 
1_1010010101010010

1_1010010101010010 + 0_1101011011111010 = 
0111110001001100

0111110001001100 >> 1 = 
0011111000100110


// ---------------------------------------------------------------------------------------------------------------------------------------



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0100101011110100
D[WIDTH-1:0] = 0000000000000010
Q[WIDTH-1:0] = X / D = 0010010101111010
REM[WIDTH-1:0] = 0000000000000000

CLZ_X = 1
CLZ_D = 14
CLZ_DIFF = CLZ_D - CLZ_X = 13
Normalized_D = 1000000000000000
根据D的值, 可得选择常数:
m[-1] = -13
m[ 0] = - 4
m[+1] = + 4
m[+2] = +12

+ D[ITN_W-1:0] = 0_1000000000000000
+2D[ITN_W-1:0] = 1_0000000000000000
- D[ITN_W-1:0] = 1_1000000000000000
-2D[ITN_W-1:0] = 1_0000000000000000
~2D[ITN_W-1:0] = 0_1111111111111111

l_shift_num = CLZ_D = 1
shifted_dividend[(2 * WIDTH + 1)-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000000100101011110100 << 14 = 
0_00010010101111010000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w[0][ITN_W-1:0] = 0_0001001010111101
(4 * w[0])_trunc_3_4 = 000_0100, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
0000000000000000

ITER[0]:
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_0100101011110100 + 
1_1000000000000000 = 
1_1100101011110100
(4 * w[1])_trunc_3_4 = 111_0010, "belongs to [-Inf, m[-1])" -> q[2] = -2
q_pos = 0100
q_neg = 0010
temp_dividend[1][WIDTH-1:0] = temp_dividend[0][WIDTH-1:0] << 2 = 
0000000000000000

ITER[1]:
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
1_0010101111010000 + 
1_0000000000000000 = 
0_0010101111010000
(4 * w[2])_trunc_3_4 = 000_1010, "belongs to [m[+1], m[+2])" -> q[3] = +1
q_pos = 0100_01
q_neg = 0010_00
temp_dividend[2][WIDTH-1:0] = temp_dividend[1][WIDTH-1:0] << 2 = 
0000000000000000

ITER[2]:
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_1010111101000000 + 
1_1000000000000000 = 
0_0010111101000000
(4 * w[3])_trunc_3_4 = 000_1011, "belongs to [m[+1], m[+2])" -> q[4] = +1
q_pos = 0100_0101
q_neg = 0010_0000
temp_dividend[3][WIDTH-1:0] = temp_dividend[2][WIDTH-1:0] << 2 = 
0000000000000000

ITER[3]:
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_1011110100000000 + 
1_1000000000000000 = 
0_0011110100000000
(4 * w[4])_trunc_3_4 = 000_1111, "belongs to [m[+2], +Inf)" -> q[5] = +2
q_pos = 0100_0101_10
q_neg = 0010_0000_00
temp_dividend[4][WIDTH-1:0] = temp_dividend[3][WIDTH-1:0] << 2 = 
0000000000000000

ITER[4]:
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_1111010000000000 + 
1_0000000000000000 = 
1_1111010000000000
(4 * w[5])_trunc_3_4 = 111_1101, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0100_0101_1000
q_neg = 0010_0000_0000
temp_dividend[5][WIDTH-1:0] = temp_dividend[4][WIDTH-1:0] << 2 = 
0000000000000000

ITER[5]:
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
1_1101000000000000 + 
0_0000000000000000 = 
1_1101000000000000
(4 * w[6])_trunc_3_4 = 111_0100, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0100_0101_1000_00
q_neg = 0010_0000_0000_01
temp_dividend[6][WIDTH-1:0] = temp_dividend[5][WIDTH-1:0] << 2 = 
0000000000000000

ITER[6]:
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
1_0100000000000000 + 
0_1000000000000000 = 
1_1100000000000000
(4 * w[7])_trunc_3_4 = 111_0000, "belongs to [-Inf, m[-1])" -> q[8] = -2
q_pos = 0100_0101_1000_0000
q_neg = 0010_0000_0000_0110
temp_dividend[7][WIDTH-1:0] = temp_dividend[6][WIDTH-1:0] << 2 = 
0000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
1_0000000000000000 + 
1_0000000000000000 = 
0_0000000000000000 >= 0

corr(q_pos - q_neg) = 0010010101111010


// ---------------------------------------------------------------------------------------------------------------------------------------















算法原理链接:
https://digitalsystemdesign.in/signed-array-divider/


// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 32;
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 10000001010111000000011000101110 = 2170291758
D[WIDTH-1:0] = 00000001001101000001100110100011 = 20191651
Q[WIDTH-1:0] = X / D = 107 = 00000000000000000000000001101011
REM[WIDTH-1:0] = 2170291758 - 20191651 * 107 = 9785101 = 00000000100101010100111100001101


stage[0]:
|(D[31:1]) = 1 -> rem[0] = X[31] = 1
q[31] = 0
q = 0

stage[1]:
{rem[0], X[30]} - D[1:0] = 
10 - 
11 = 
1_11 < 0, |(D[31:2]) = 1
rem[1] = 10
q[30] = 0
q = 00

stage[2]:
{rem[1], X[29]} - D[2:0] = 
100 - 
011 = 
0_001 >= 0, |(D[31:3]) = 1
rem[2] = 100
q[29] = 0
q = 000

stage[3]:
{rem[2], X[28]} - D[3:0] = 
1000 - 
0011 = 
0_0101 >= 0, |(D[31:4]) = 1
rem[3] = 1000
q[28] = 0
q = 0000

stage[4]:
{rem[3], X[27]} - D[4:0] = 
10000 - 
00011 = 
0_01101 >= 0, |(D[31:5]) = 1
rem[4] = 10000
q[27] = 0
q = 0000_0

stage[5]:
{rem[4], X[26]} - D[5:0] = 
100000 - 
100011 = 
1_111101 < 0, |(D[31:6]) = 1
rem[5] = 100000
q[26] = 0
q = 0000_00

stage[6]:
{rem[5], X[25]} - D[6:0] = 
1000000 - 
0100011 = 
0_0011101 >= 0, |(D[31:7]) = 1
rem[6] = 1000000
q[25] = 0
q = 0000_000

stage[7]:
{rem[6], X[24]} - D[7:0] = 
10000001 - 
10100011 = 
1_11011110 < 0, |(D[31:8]) = 1
rem[7] = 10000001
q[24] = 0
q = 0000_0000

stage[8]:
{rem[7], X[23]} - D[8:0] = 
100000010 - 
110100011 = 
1_101011111 < 0, |(D[31:9]) = 1
rem[8] = 100000010
q[23] = 0
q = 0000_0000_0

stage[9]:
{rem[8], X[22]} - D[9:0] = 
1000000101 - 
0110100011 = 
0_0001100010 >= 0, |(D[31:10]) = 1
rem[9] = 1000000101
q[22] = 0
q = 0000_0000_00

stage[10]:
{rem[9], X[21]} - D[10:0] = 
10000001010 - 
00110100011 = 
0_01001100111 >= 0, |(D[31:11]) = 1
rem[10] = 10000001010
q[21] = 0
q = 0000_0000_000

stage[11]:
{rem[10], X[20]} - D[11:0] = 
100000010101 - 
100110100011 = 
1_111001110010 < 0, |(D[31:12]) = 1
rem[11] = 100000010101
q[20] = 0
q = 0000_0000_0000

stage[12]:
{rem[11], X[19]} - D[12:0] = 
1000000101011 - 
1100110100011 = 
1_1011010001000 < 0, |(D[31:13]) = 1
rem[12] = 1000000101011
q[19] = 0
q = 0000_0000_0000_0

stage[13]:
{rem[12], X[18]} - D[13:0] = 
10000001010111 - 
01100110100011 = 
0_00011010110100 >= 0, |(D[31:14]) = 1
rem[13] = 10000001010111
q[18] = 0
q = 0000_0000_0000_00

stage[14]:
{rem[13], X[17]} - D[14:0] = 
100000010101110 - 
001100110100011 = 
0_010011100001011 >= 0, |(D[31:15]) = 1
rem[14] = 100000010101110
q[17] = 0
q = 0000_0000_0000_000

stage[15]:
{rem[14], X[16]} - D[15:0] = 
1000000101011100 - 
0001100110100011 = 
0_0110011110111001 >= 0, |(D[31:16]) = 1
rem[15] = 1000000101011100
q[16] = 0
q = 0000_0000_0000_0000

stage[16]:
{rem[15], X[15]} - D[16:0] = 
10000001010111000 - 
00001100110100011 = 
0_01110100100010101 >= 0, |(D[31:17]) = 1
rem[16] = 10000001010111000
q[15] = 0
q = 0000_0000_0000_0000_0

stage[17]:
{rem[16], X[14]} - D[17:0] = 
100000010101110000 - 
000001100110100011 = 
0_011110101111001101 >= 0, |(D[31:18]) = 1
rem[17] = 100000010101110000
q[14] = 0
q = 0000_0000_0000_0000_00

stage[18]:
{rem[17], X[13]} - D[18:0] = 
1000000101011100000 - 
1000001100110100011 = 
1_1111111000100111101 < 0, |(D[31:19]) = 1
rem[18] = 1000000101011100000
q[13] = 0
q = 0000_0000_0000_0000_000

stage[19]:
{rem[18], X[12]} - D[19:0] = 
10000001010111000000 - 
01000001100110100011 = 
0_00111111110000011101 >= 0, |(D[31:20]) = 1
rem[20] = 10000001010111000000
q[12] = 0
q = 0000_0000_0000_0000_0000

stage[20]:
{rem[19], X[11]} - D[20:0] = 
100000010101110000000 - 
101000001100110100011 = 
1_111000001000111011101 < 0, |(D[31:21]) = 1
rem[20] = 100000010101110000000
q[11] = 0
q = 0000_0000_0000_0000_0000_0

stage[21]:
{rem[20], X[10]} - D[21:0] = 
1000000101011100000001 - 
1101000001100110100011 = 
1_1011000011110101011110 < 0, |(D[31:22]) = 1
rem[21] = 1000000101011100000001
q[10] = 0
q = 0000_0000_0000_0000_0000_00

stage[22]:
{rem[21], X[9]} - D[22:0] = 
10000001010111000000011 - 
01101000001100110100011 = 
0_00011001001010001100000 >= 0, |(D[31:23]) = 1
rem[22] = 10000001010111000000011
q[9] = 0
q = 0000_0000_0000_0000_0000_000

stage[23]:
{rem[22], X[8]} - D[23:0] = 
100000010101110000000110 - 
001101000001100110100011 = 
0_010011010100001001100011 >= 0, |(D[31:24]) = 1
rem[23] = 100000010101110000000110
q[8] = 0
q = 0000_0000_0000_0000_0000_0000

stage[24]:
{rem[23], X[7]} - D[24:0] = 
1000000101011100000001100 - 
1001101000001100110100011 = 
1_1110011101001111001101001 < 0, |(D[31:25]) = 0
rem[24] = 1000000101011100000001100
q[7] = 0
q = 0000_0000_0000_0000_0000_0000_0

stage[25]:
{rem[24], X[6]} - D[25:0] = 
10000001010111000000011000 - 
01001101000001100110100011 = 
0_00110100010101011001110101 >= 0, |(D[31:26]) = 0
rem[25] = 00110100010101011001110101
q[6] = 1
q = 0000_0000_0000_0000_0000_0000_01

stage[26]:
{rem[25], X[5]} - D[26:0] = 
001101000101010110011101011 - 
001001101000001100110100011 = 
0_000011011101001001101001000 >= 0, |(D[31:27]) = 0
rem[26] = 000011011101001001101001000
q[5] = 1
q = 0000_0000_0000_0000_0000_0000_011

stage[27]:
{rem[26], X[4]} - D[27:0] = 
0000110111010010011010010000 - 
0001001101000001100110100011 = 
1_1111101010010000110011101101 < 0, |(D[31:28]) = 0
rem[27] = 0000110111010010011010010000
q[4] = 0
q = 0000_0000_0000_0000_0000_0000_0110

stage[28]:
{rem[27], X[3]} - D[28:0] = 
00001101110100100110100100001 - 
00001001101000001100110100011 = 
0_00000100001100011001101111110 >= 0, |(D[31:29]) = 0
rem[28] = 00000100001100011001101111110
q[3] = 1
q = 0000_0000_0000_0000_0000_0000_0110_1

stage[29]:
{rem[28], X[2]} - D[29:0] = 
000001000011000110011011111101 - 
000001001101000001100110100011 = 
1_111111110110000100110101011010 < 0, |(D[31:30]) = 0
rem[29] = 000001000011000110011011111101
q[2] = 0
q = 0000_0000_0000_0000_0000_0000_0110_10

stage[30]:
{rem[29], X[1]} - D[30:0] = 
0000010000110001100110111111011 - 
0000001001101000001100110100011 = 
0_0000000111001001011010001011000 >= 0, |(D[31:31]) = 0
rem[30] = 0000000111001001011010001011000
q[1] = 1
q = 0000_0000_0000_0000_0000_0000_0110_101

stage[31]:
{rem[30], X[0]} - D[30:0] = 
00000001110010010110100010110000 - 
00000001001101000001100110100011 = 
0_00000000100101010100111100001101 >= 0
rem[31] = 00000000100101010100111100001101
q[0] = 1
q = 0000_0000_0000_0000_0000_0000_0110_1011

q_final = 00000000000000000000000001101011

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 10001101010111000110011010001001 = 2371643017
D[WIDTH-1:0] = 00000000000000000000000000000011 = 3
Q[WIDTH-1:0] = X / D = 790547672 = 00101111000111101100110011011000
REM[WIDTH-1:0] = 2371643017 - 790547672 * 3 = 1 = 00000000000000000000000000000001


stage[0]:
|(D[31:1]) = 1 -> rem[0] = X[31] = 1
q = 0

stage[1]:
{rem[0], X[30]} - D[1:0] = 
10 - 
11 = 
1_11 < 0, |(D[31:2]) = 0
rem[1] = 10
q = 00

stage[2]:
{rem[1], X[29]} - D[2:0] = 
100 - 
011 = 
0_001 >= 0, |(D[31:3]) = 0
rem[2] = 001
q = 001

stage[3]:
{rem[2], X[28]} - D[3:0] = 
0010 - 
0011 = 
1_1111 < 0, |(D[31:4]) = 0
rem[3] = 0010
q = 0010

stage[4]:
{rem[3], X[27]} - D[4:0] = 
00101 - 
00011 = 
0_00010 >= 0, |(D[31:5]) = 0
rem[4] = 00010
q = 00101

stage[5]:
{rem[4], X[26]} - D[5:0] = 
000101 - 
000011 = 
0_000010 >= 0, |(D[31:6]) = 0
rem[5] = 000010
q = 001011

stage[6]:
{rem[5], X[25]} - D[6:0] = 
0000100 - 
0000011 = 
0_0000001 >= 0, |(D[31:7]) = 0
rem[6] = 0000001
q = 0010111

stage[7]:
{rem[6], X[24]} - D[7:0] = 
00000011 - 
00000011 = 
0_00000000 >= 0, |(D[31:8]) = 0
rem[7] = 00000000
q = 00101111

stage[8]:
{rem[7], X[23]} - D[8:0] = 
000000000 - 
000000011 = 
1_111111101 < 0, |(D[31:9]) = 0
rem[8] = 000000000
q = 001011110

stage[9]:
{rem[8], X[22]} - D[9:0] = 
0000000001 - 
0000000011 = 
1_1111111110 < 0, |(D[31:10]) = 0
rem[9] = 0000000001
q = 0010111100

stage[10]:
{rem[9], X[21]} - D[10:0] = 
00000000010 - 
00000000011 = 
1_11111111111 < 0, |(D[31:11]) = 0
rem[10] = 00000000010
q = 00101111000

stage[11]:
{rem[10], X[20]} - D[11:0] = 
000000000101 - 
000000000011 = 
0_000000000010 >= 0, |(D[31:12]) = 0
rem[11] = 000000000010
q = 001011110001

stage[12]:
{rem[11], X[19]} - D[12:0] = 
0000000000101 - 
0000000000011 = 
0_0000000000010 >= 0, |(D[31:13]) = 0
rem[12] = 0000000000010
q = 0010111100011

stage[13]:
{rem[12], X[18]} - D[13:0] = 
00000000000101 - 
00000000000011 = 
0_00000000000010 >= 0, |(D[31:14]) = 0
rem[13] = 00000000000010
q = 00101111000111

stage[14]:
{rem[13], X[17]} - D[14:0] = 
000000000000100 - 
000000000000011 = 
0_000000000000001 >= 0, |(D[31:15]) = 0
rem[14] = 000000000000001
q = 001011110001111

stage[15]:
{rem[14], X[16]} - D[15:0] = 
0000000000000010 - 
0000000000000011 = 
1_1111111111111111 < 0, |(D[31:16]) = 0
rem[15] = 0000000000000010
q = 0010111100011110

stage[16]:
{rem[15], X[15]} - D[16:0] = 
00000000000000100 - 
00000000000000011 = 
0_00000000000000001 >= 0, |(D[31:17]) = 0
rem[16] = 00000000000000001
q = 00101111000111101

stage[17]:
{rem[16], X[14]} - D[17:0] = 
000000000000000011 - 
000000000000000011 = 
0_000000000000000000 >= 0, |(D[31:18]) = 0
rem[17] = 000000000000000000
q = 001011110001111011

stage[18]:
{rem[17], X[13]} - D[18:0] = 
0000000000000000001 - 
0000000000000000011 = 
1_1111111111111111110 < 0, |(D[31:19]) = 0
rem[18] = 0000000000000000001
q = 0010111100011110110

stage[19]:
{rem[18], X[12]} - D[19:0] = 
00000000000000000010 - 
00000000000000000011 = 
1_11111111111111111111 < 0, |(D[31:20]) = 0
rem[20] = 00000000000000000010
q = 00101111000111101100

stage[20]:
{rem[19], X[11]} - D[20:0] = 
000000000000000000100 - 
000000000000000000011 = 
0_000000000000000000001 >= 0, |(D[31:21]) = 0
rem[20] = 000000000000000000001
q = 001011110001111011001

stage[21]:
{rem[20], X[10]} - D[21:0] = 
0000000000000000000011 - 
0000000000000000000011 = 
0_0000000000000000000000 >= 0 |(D[31:22]) = 0
rem[21] = 0000000000000000000000
q = 0010111100011110110011

stage[22]:
{rem[21], X[9]} - D[22:0] = 
00000000000000000000001 - 
00000000000000000000011 = 
1_11111111111111111111110 < 0, |(D[31:23]) = 0
rem[22] = 00000000000000000000001
q = 00101111000111101100110

stage[23]:
{rem[22], X[8]} - D[23:0] = 
000000000000000000000010 - 
000000000000000000000011 = 
1_111111111111111111111111 < 0, |(D[31:24]) = 0
rem[23] = 000000000000000000000010
q = 001011110001111011001100

stage[24]:
{rem[23], X[7]} - D[24:0] = 
0000000000000000000000101 - 
0000000000000000000000011 = 
0_0000000000000000000000010 >= 0, |(D[31:25]) = 0
rem[24] = 0000000000000000000000010
q = 0010111100011110110011001

stage[25]:
{rem[24], X[6]} - D[25:0] = 
00000000000000000000000100 - 
00000000000000000000000011 = 
0_00000000000000000000000001 >= 0, |(D[31:26]) = 0
rem[25] = 00000000000000000000000001
q = 00101111000111101100110011

stage[26]:
{rem[25], X[5]} - D[26:0] = 
000000000000000000000000010 - 
000000000000000000000000011 = 
1_111111111111111111111111111 < 0, |(D[31:27]) = 0
rem[26] = 000000000000000000000000010
q = 001011110001111011001100110

stage[27]:
{rem[26], X[4]} - D[27:0] = 
0000000000000000000000000100 - 
0000000000000000000000000011 = 
0_0000000000000000000000000001 >= 0, |(D[31:28]) = 0
rem[27] = 0000000000000000000000000001
q = 0010111100011110110011001101

stage[28]:
{rem[27], X[3]} - D[28:0] = 
00000000000000000000000000011 - 
00000000000000000000000000011 = 
0_00000000000000000000000000000 >= 0, |(D[31:29]) = 0
rem[28] = 00000000000000000000000000000
q = 00101111000111101100110011011

stage[29]:
{rem[28], X[2]} - D[29:0] = 
000000000000000000000000000000 - 
000000000000000000000000000011 = 
1_111111111111111111111111111101 < 0, |(D[31:30]) = 0
rem[29] = 000000000000000000000000000000
q = 001011110001111011001100110110

stage[30]:
{rem[29], X[1]} - D[30:0] = 
0000000000000000000000000000000 - 
0000000000000000000000000000011 = 
1_1111111111111111111111111111101 < 0, |(D[31:31]) = 0
rem[30] = 0000000000000000000000000000000
q = 0010111100011110110011001101100

stage[31]:
{rem[30], X[0]} - D[30:0] = 
00000000000000000000000000000001 - 
00000000000000000000000000000011 = 
1_11111111111111111111111111111110 < 0
rem[31] = 00000000000000000000000000000001
q = 00101111000111101100110011011000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 11111101011111000110011011110011 = 4252788467
D[WIDTH-1:0] = 00000000000000000010011001001001 = 9801
Q[WIDTH-1:0] = X / D = 433913 = 00000000000001101001111011111001
REM[WIDTH-1:0] = 4252788467 - 9801 * 433913 = 7154 = 00000000000000000001101111110010

stage[0]:
|(D[31:1]) = 1 -> rem[0] = X[31] = 1
q = 0

stage[1]:
{rem[0], X[30]} - D[1:0] = 
11 - 
01 = 
0_10 >= 0, |(D[31:2]) = 1
rem[1] = 11
q = 00

stage[2]:
{rem[1], X[29]} - D[2:0] = 
111 - 
001 = 
0_110 >= 0, |(D[31:3]) = 1
rem[2] = 111
q = 000

stage[3]:
{rem[2], X[28]} - D[3:0] = 
1111 - 
1001 = 
0_0110 >= 0, |(D[31:4]) = 1
rem[3] = 1111
q = 0000

stage[4]:
{rem[3], X[27]} - D[4:0] = 
11111 - 
01001 = 
0_10110 >= 0, |(D[31:5]) = 1
rem[4] = 11111
q = 00000

stage[5]:
{rem[4], X[26]} - D[5:0] = 
111111 - 
001001 = 
0_110110 >= 0, |(D[31:6]) = 1
rem[5] = 111111
q = 000000

stage[6]:
{rem[5], X[25]} - D[6:0] = 
1111110 - 
1001001 = 
0_01101011 >= 0, |(D[31:7]) = 1
rem[6] = 1111110
q = 0000000

stage[7]:
{rem[6], X[24]} - D[7:0] = 
11111101 - 
01001001 = 
0_10110100 >= 0, |(D[31:8]) = 1
rem[7] = 11111101
q = 00000000

stage[8]:
{rem[7], X[23]} - D[8:0] = 
111111010 - 
001001001 = 
0_110110001 >= 0, |(D[31:9]) = 1
rem[8] = 111111010
q = 000000000

stage[9]:
{rem[8], X[22]} - D[9:0] = 
1111110101 - 
1001001001 = 
0_0110101100 >= 0, |(D[31:10]) = 1
rem[9] = 1111110101
q = 0000000000

stage[10]:
{rem[9], X[21]} - D[10:0] = 
11111101011 - 
11001001001 = 
0_00110100010 >= 0, |(D[31:11]) = 1
rem[10] = 11111101011
q = 00000000000

stage[11]:
{rem[10], X[20]} - D[11:0] = 
111111010111 - 
011001001001 = 
0_100110001110 >= 0, |(D[31:12]) = 1
rem[11] = 111111010111
q = 000000000000

stage[12]:
{rem[11], X[19]} - D[12:0] = 
1111110101111 - 
0011001001001 = 
0_1100101100110 >= 0, |(D[31:13]) = 1
rem[12] = 1111110101111
q = 0000000000000

stage[13]:
{rem[12], X[18]} - D[13:0] = 
11111101011111 - 
10011001001001 = 
0_01100100010110 >= 0, |(D[31:14]) = 0
rem[13] = 01100100010110
q = 00000000000001

stage[14]:
{rem[13], X[17]} - D[14:0] = 
011001000101100 - 
010011001001001 = 
0_000101111100011 >= 0, |(D[31:15]) = 0
rem[14] = 000101111100011
q = 000000000000011

stage[15]:
{rem[14], X[16]} - D[15:0] = 
0001011111000110 - 
0010011001001001 = 
1_1111000101111101 < 0, |(D[31:16]) = 0
rem[15] = 0001011111000110
q = 0000000000000110

stage[16]:
{rem[15], X[15]} - D[16:0] = 
00010111110001100 - 
00010011001001001 = 
0_00000100101000011 >= 0, |(D[31:17]) = 0
rem[16] = 00000100101000011
q = 00000000000001101

stage[17]:
{rem[16], X[14]} - D[17:0] = 
000001001010000111 - 
000010011001001001 = 
1_111110110000111110 < 0, |(D[31:18]) = 0
rem[17] = 000001001010000111
q = 000000000000011010

stage[18]:
{rem[17], X[13]} - D[18:0] = 
0000010010100001111 - 
0000010011001001001 = 
1_1111111111011000110 < 0, |(D[31:19]) = 0
rem[18] = 0000010010100001111
q = 0000000000000110100

stage[19]:
{rem[18], X[12]} - D[19:0] = 
00000100101000011110 - 
00000010011001001001 = 
0_00000010001111010101 >= 0, |(D[31:20]) = 0
rem[20] = 00000010001111010101
q = 00000000000001101001

stage[20]:
{rem[19], X[11]} - D[20:0] = 
000000100011110101010 - 
000000010011001001001 = 
0_000000010000101100001 >= 0, |(D[31:21]) = 0
rem[20] = 000000010000101100001
q = 000000000000011010011

stage[21]:
{rem[20], X[10]} - D[21:0] = 
0000000100001011000011 - 
0000000010011001001001 = 
0_0000000001110001111010 >= 0 |(D[31:22]) = 0
rem[21] = 0000000001110001111010
q = 0000000000000110100111

stage[22]:
{rem[21], X[9]} - D[22:0] = 
00000000011100011110101 - 
00000000010011001001001 = 
0_00000000001001010101100 >= 0, |(D[31:23]) = 0
rem[22] = 00000000001001010101100
q = 00000000000001101001111

stage[23]:
{rem[22], X[8]} - D[23:0] = 
000000000010010101011000 - 
000000000010011001001001 = 
1_111111111111111100001111 < 0, |(D[31:24]) = 0
rem[23] = 000000000010010101011000
q = 000000000000011010011110

stage[24]:
{rem[23], X[7]} - D[24:0] = 
0000000000100101010110001 - 
0000000000010011001001001 = 
0_0000000000010010001101000 >= 0, |(D[31:25]) = 0
rem[24] = 0000000000010010001101000
q = 0000000000000110100111101

stage[25]:
{rem[24], X[6]} - D[25:0] = 
00000000000100100011010001 - 
00000000000010011001001001 = 
0_00000000000010001010001000 >= 0, |(D[31:26]) = 0
rem[25] = 00000000000010001010001000
q = 00000000000001101001111011

stage[26]:
{rem[25], X[5]} - D[26:0] = 
000000000000100010100010001 - 
000000000000010011001001001 = 
0_000000000000001111011001000 >= 0, |(D[31:27]) = 0
rem[26] = 000000000000001111011001000
q = 000000000000011010011110111

stage[27]:
{rem[26], X[4]} - D[27:0] = 
0000000000000011110110010001 - 
0000000000000010011001001001 = 
0_0000000000000001011101001000 >= 0, |(D[31:28]) = 0
rem[27] = 0000000000000001011101001000
q = 0000000000000110100111101111

stage[28]:
{rem[27], X[3]} - D[28:0] = 
00000000000000010111010010000 - 
00000000000000010011001001001 = 
0_00000000000000000100001000111 >= 0, |(D[31:29]) = 0
rem[28] = 00000000000000000100001000111
q = 00000000000001101001111011111

stage[29]:
{rem[28], X[2]} - D[29:0] = 
000000000000000001000010001110 - 
000000000000000010011001001001 = 
1_111111111111111110101001000101 < 0, |(D[31:30]) = 0
rem[29] = 000000000000000001000010001110
q = 000000000000011010011110111110

stage[30]:
{rem[29], X[1]} - D[30:0] = 
0000000000000000010000100011101 - 
0000000000000000010011001001001 = 
1_1111111111111111111101011010100 < 0, |(D[31:31]) = 0
rem[30] = 0000000000000000010000100011101
q = 0000000000000110100111101111100

stage[31]:
{rem[30], X[0]} - D[30:0] = 
00000000000000000100001000111011 - 
00000000000000000010011001001001 = 
0_00000000000000000001101111110010 >= 0
rem[31] = 00000000000000000001101111110010
q = 00000000000001101001111011111001



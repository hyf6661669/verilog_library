

a0[3:0] = 11 = 1011
b0[3:0] = 5 = 0101
a1[3:0] = 8 = 1000
b1[3:0] = 5 = 0101
a2[3:0] = 3 = 0011
b2[3:0] = 9 = 1001
a3[3:0] = 12 = 1100
b3[3:0] = 4 = 0100

有以下属性:
(a0 + b0) == 0
(a1 + b1) != 0
(a2 + b2) != 0
(a3 + b3) == 0

a_merged[15:0] = {a3, a2, a1, a0} = 1100001110001011
b_merged[15:0] = {a3, a2, a1, a0} = 0100100101010101

a_merged[15:1] ^ b_merged[15:1] = 100010101101111
a_merged[14:0] | b_merged[14:0] = 100101111011111

a[15:0] = 65530 = 1111111111111010
b[15:0] = 6 = 0000000000000110

a[15:1] ^ b[15:1] = 111111111111110
a[15:1] | b[15:1] = 111111111111110

对于I16的数据来说, 需要检查XOR/OR结果的[14:0], 那么才能知道((ax + bx) == 0)的结果


a0[3:0] = 11 = 1011
b0[3:0] = 5 = 0101
a1[3:0] = 7 = 0111
b1[3:0] = 9 = 1001
a2[3:0] = 3 = 0011
b2[3:0] = 13 = 1101
a3[3:0] = 12 = 1100
b3[3:0] = 4 = 0100

a_merged[15:0] = {a3, a2, a1, a0} = 1100001101111011
b_merged[15:0] = {b3, b2, b1, b0} = 0100110110010101

a_merged[15:1] ^ b_merged[15:1] = 100_0_111_0_111_0_111
a_merged[14:0] | b_merged[14:0] = 100_1_111_1_111_1_111

对于I4的数据来说, 如果只检查XOR/OR结果的[14:12], [10:8], [6:4], [2:0], 那么才能知道((ax + bx) == 0)的结果

假设有2个11-bit的I11数据和4个I4数据共用一个XOR/OR逻辑:
a[10:0] = 1055 = 10000011111
b[10:0] = 2048 - 1055 = 983 = 01111100001

a_merged[15:0] = {a[10:0], 5'b0} = 1000001111100000
b_merged[15:0] = {b[10:0], 5'b0} = 0111110000100000

a_merged[15:1] ^ b_merged[15:1] = 111_1_111_1_110_0_000
a_merged[14:0] | b_merged[14:0] = 111_1_111_1_110_0_000



// 综上所述应当将XOR/OR结果分为5部分, 根据fp_fmt的值来决定使用哪些部分

// a_merged_v2[18:0] = {a3, 0, a2, 0, a1, 0, a0} = 1100_0_0011_0_0111_0_1011
// b_merged_v2[18:0] = {b3, 0, b2, 0, b1, 0, b0} = 0100_0_1101_0_1001_0_0101

// a_merged_v2[18:1] ^ a_merged_v2[18:1] = 100001110011100111
// a_merged_v2[17:0] | a_merged_v2[17:0] = 100011110111101111

// ================================================================================================================================================
// ================================================================================================================================================
// ================================================================================================================================================
// ================================================================================================================================================
93.4ns
121.6ns
// ================================================================================================================================================

ref_res = 20782081 = 0_01000000_11110000010000010000001

rt_q = f8208208b9d178 = 11111000001000001000001000_001000101110011101000101111000


rt_m1_q = 1e082070b9d174 = 1111000001000001000000111_0000101110011101000101110100







rt_m1_pre_inc_0 = c8f1508b73464 = 110010001111000101010000_1_000101101110011010001100100



sum = ca6e97b052e610f0 = 1100101001101110100101111011_000001010010111001100001000011110000
cry = 372a80109ae38c80 = 0011011100101010100000000001_000010011010111000111000110010000000

1100101001101110100101111011 + 
0011011100101010100000000001 = 
0000000110011001000101111100

ref_sum = c66ee840003fff = 11000110011011101110100001000000000000000011111111111111
ref_cry = 372a2f7fffc001 = 00110111001010100010111101111111111111111100000000000001



ref_frac = 1.11001000111100010101000_0111111010100111100000000


cyc[0]: 
f_r_s_for_csa_0[1] = 07f00004c23f80 = 0000011111110000000000000000_0100110000100011111110000000
f_r_c_for_csa_0[1] = 0000000c000000 = 0000000000000000000000000000_1100000000000000000000000000

sqrt_csa_val[0] = f0000010000000 = 1111000000000000000000000001_0000000000000000000000000000



dut_sum = f08dafb0 = 11110000100011011010111110110000
dut_cry = 1ce4a090 = 00011100111001001010000010010000
addend = 00001101011100100101000001000000

ref_sum = f08dafffffffff = 11110000100011011010111111111111111111111111111111111111
ref_cry = 1ce4a000000001 = 00011100111001001010000000000000000000000000000000000001
addend = 00001101011100100101000000000000000000000000000000000000

a_frac = 10101001100101010101010101001100101010101010101001100
sqrt(a_frac) = 1.0010011010101001111001001111000011100000000001101000_101001001110110001010101...

init_rem_sum_noadj = 000010100110010101010101010100110010101010101010100110000000000

// ================================================================================================================================================
// iter[0]:
// ================================================================================================================================================
rem_sum_f3 = 000010100110010101010101010100110010101010101010100110000000000
rem_carry_f3 = 000000000000000000000000000000000000000000000000000000000000000

raw_mask_f3 = 000000000000000000
quot_f3 = 1000000000000000000000000000000000000000000000000000000
quot_m1_f3 = 0000000000000000000000000000000000000000000000000000000

mask_f3[0] = 10000000000000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
10000000000000000000000000000000000000000000000000000000 ^ 
11000000000000000000000000000000000000000000000000000000 = 
01000000000000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0100000000000000000000000000000000000000000000000000000 |
1000000000000000000000000000000000000000000000000000000 = 
1100000000000000000000000000000000000000000000000000000

mask_f3[1] 		= 11000000000000000000000000000000000000000000000000000000
msk_dig[1] 		= 00100000000000000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0110000000000000000000000000000000000000000000000000000

mask_f3[2] 		= 11100000000000000000000000000000000000000000000000000000
msk_dig[2] 		= 00010000000000000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0011000000000000000000000000000000000000000000000000000


rem_sum_f3[62:60] = 000
rem_carry_f3[62:60] = 000
-> 
quot_dig0[0] = 01
->
prev_quot[0] = quot_f3 = 1000000000000000000000000000000000000000000000000000000
prev_quot_m1[0] = quot_m1_f3 = 0000000000000000000000000000000000000000000000000000000
new_quot0_f3[0] = prev_quot[0] & mask_f3[0][55:1] | msk_dig[0][55:1] = 1100000000000000000000000000000000000000000000000000000
new_quot0_m1_f3[0] = prev_quot[0] & mask_f3[0][55:1] = 1000000000000000000000000000000000000000000000000000000

csa_minus_val_sqrt0[0] = {quot_f3[53: 1], 2'b0} | msk_dig[0][55: 1] = 
0000000000000000000000000000000000000000000000000000000 | 
0100000000000000000000000000000000000000000000000000000 = 
0100000000000000000000000000000000000000000000000000000
csa_val0[0] = ~csa_minus_val0[0][50:0] = 111111111111111111111111111111111111111111111111111
csa_mux[0] = 111111111111111111111111111111111111111111111111111000000

rem_sum_in[0] = rem_sum_f3[61:0] = 00010100110010101010101010100110010101010101010100110000000000
rem_carry_in[0] = rem_carry_f3[61:0] = 00000000000000000000000000000000000000000000000000000000000000

rem_sum_in[0][61:56] 		= 000101
rem_carry_in[0][61:56] 		= 000000
csa_minus_val0[0][54:51] 	=   0100 -> 1011
rem0_sum_minus[0][5:0] 		= 001110
rem0_carry_minus[0][5:0] 	= 100011
rem_sum_msb0[0][5:0] 		= 001110
rem_carry_msb0[0][5:0] 		= 100011


rem_sum_xor[0][56:0] = 
001100101010101010101001100101010101010101001100000000000 ^ 
000000000000000000000000000000000000000000000000000000000 ^ 
111111111111111111111111111111111111111111111111111000000 = 
110011010101010101010110011010101010101010110011111000000
rem_carry_andor[0][57:0] = 0011001010101010101010011001010101010101010011000000000001


new_rem_sum0[0][56:0] = {rem_sum_msb0[0][5:0], rem_sum_xor[0][56: 6]} = 001110110011010101010101010110011010101010101010110011111
new_rem_sum_f3[0] = {new_rem_sum0[0][56:0], 6'b0} = 001110110011010101010101010110011010101010101010110011111000000
new_rem_carry0[0][55:0] = {rem_carry_msb0[0][5:1], rem_carry_andor[0][57: 7]} = 10001001100101010101010101001100101010101010101001100000
new_rem_carry_f3[0] = {new_rem_carry0[0][55:0], quot_dig0[0][0], 6'b0} = 100010011001010101010101010011001010101010101010011000001000000


new_rem_sum_f3[0] + new_rem_carry_f3[0] = 
001110110011010101010101010110011010101010101010110011111000000 + 
100010011001010101010101010011001010101010101010011000001000000 = 
110001001100101010101010101001100101010101010101001100000000000
{1'b0, ({new_quot0_m1_f3[0], 1'b0} | msk_dig[1]), 6'b0} = 010100000000000000000000000000000000000000000000000000000000000

110001001100101010101010101001100101010101010101001100000000000 + 
010100000000000000000000000000000000000000000000000000000000000 = 
000101001100101010101010101001100101010101010101001100000000000
000101001100101010101010101001100101010101010101001100

// ====================================
rem_sum_in[1] = new_rem_sum_f3[0][61:0] = 01110110011010101010101010110011010101010101010110011111000000
rem_carry_in[1] = new_rem_carry_f3[0][61:0] = 00010011001010101010101010011001010101010101010011000001000000

rem_sum_msb0[0][5:3] = 001
rem_carry_msb0[0][5:3] = 100
->
quot_dig0[1] = 10
->
prev_quot[1] = new_quot0_f3[0] = 1100000000000000000000000000000000000000000000000000000
prev_quot_m1[1] = new_quot0_m1_f3[0] = 1000000000000000000000000000000000000000000000000000000
new_quot0_f3[1] = prev_quot_m1[1] & mask_f3[1][55:1] | msk_dig[1][55:1] = 1010000000000000000000000000000000000000000000000000000
new_quot0_m1_f3[1] = prev_quot_m1[1] & mask_f3[1][55:1] = 1000000000000000000000000000000000000000000000000000000


csa_plus_val_sqrt0[1] = {new_quot0_m1_f3[0][53:1], 2'b0} | msk_dig_3[1][54: 0] = 
0000000000000000000000000000000000000000000000000000000 | 
0110000000000000000000000000000000000000000000000000000 = 
0110000000000000000000000000000000000000000000000000000
csa_val0[1] = csa_plus_val0[1][50:0] = 000000000000000000000000000000000000000000000000000
csa_mux[1] = 000000000000000000000000000000000000000000000000000000000

rem_sum_in[1][61:56] 		= 011101
rem_carry_in[1][61:56] 		= 000100
csa_plus_val0[1][54:51] 	=   0110
rem0_sum_plus[1][5:0] 		= 001111
rem0_carry_plus[1][5:0] 	= 101000
rem_sum_msb0[1][5:0] 		= 001111
rem_carry_msb0[1][5:0] 		= 101000


rem_sum_xor[1][56:0] = 
100110101010101010101100110101010101010101100111110000000 ^ 
110010101010101010100110010101010101010100110000010000000 ^ 
000000000000000000000000000000000000000000000000000000000 = 
010100000000000000001010100000000000000001010111100000000
rem_carry_andor[1][57:0] = 1000101010101010101001000101010101010101001000000100000000

new_rem_sum0[1][56:0] = {rem_sum_msb0[1][5:0], rem_sum_xor[1][56: 6]} = 001111010100000000000000001010100000000000000001010111100
new_rem_sum_f3[1] = {new_rem_sum0[1][56:0], 6'b0} = 001111010100000000000000001010100000000000000001010111100000000
new_rem_carry0[1][55:0] = {rem_carry_msb0[1][5:1], rem_carry_andor[1][57: 7]} = 10100100010101010101010100100010101010101010100100000010
new_rem_carry_f3[1] = {new_rem_carry0[1][55:0], quot_dig0[1][0], 6'b0} = 101001000101010101010101001000101010101010101001000000100000000

// ====================================
rem_sum_in[2] = new_rem_sum_f3[1][61:0] = 01111010100000000000000001010100000000000000001010111100000000
rem_carry_in[2] = new_rem_carry_f3[1][61:0] = 01001000101010101010101001000101010101010101001000000100000000

rem_sum_msb0[1][5:3] = 001
rem_carry_msb0[1][5:3] = 101
->
quot_dig0[2] = 10
->
prev_quot[2] = new_quot0_f3[1] = 1010000000000000000000000000000000000000000000000000000
prev_quot_m1[2] = new_quot0_m1_f3[1] = 1000000000000000000000000000000000000000000000000000000
new_quot0_f3[2] = prev_quot_m1[2] & mask_f3[2][55:1] | msk_dig[2][55:1] = 1001000000000000000000000000000000000000000000000000000
new_quot0_m1_f3[2] = prev_quot_m1[2] & mask_f3[2][55:1] = 1000000000000000000000000000000000000000000000000000000

csa_plus_val_sqrt0[2] = {new_quot0_m1_f3[1][53:1], 2'b0} | msk_dig_3[2][54: 0] = 
0000000000000000000000000000000000000000000000000000000 |
0011000000000000000000000000000000000000000000000000000 = 
0011000000000000000000000000000000000000000000000000000

csa_val0[2] = csa_plus_val0[2][50:0] = 000000000000000000000000000000000000000000000000000
csa_mux[1] = 000000000000000000000000000000000000000000000000000000000

rem_sum_in[2][61:56] 		= 011110
rem_carry_in[2][61:56] 		= 010010
csa_plus_val0[2][54:51] 	=   0011
rem0_sum_plus[2][5:0] 		= 011111
rem0_carry_plus[2][5:0] 	= 100100
rem_sum_msb0[2][5:0] 		= 011111
rem_carry_msb0[2][5:0] 		= 100100

rem_sum_xor[2][56:0] = 
101000000000000000010101000000000000000010101111000000000 ^ 
001010101010101010010001010101010101010010000001000000000 ^ 
000000000000000000000000000000000000000000000000000000000 = 
100010101010101010000100010101010101010000101110000000000
rem_carry_andor[2][57:0] = 0010000000000000000100010000000000000000100000010000000000

new_rem_sum0[2][56:0] = {rem_sum_msb0[2][5:0], rem_sum_xor[2][56: 6]} = 011111100010101010101010000100010101010101010000101110000
new_rem_sum_f3[2] = {new_rem_sum0[2][56:0], 6'b0} = 011111100010101010101010000100010101010101010000101110000000000
new_rem_carry0[2][55:0] = {rem_carry_msb0[2][5:1], rem_carry_andor[2][57: 7]} = 10010001000000000000000010001000000000000000010000001000
new_rem_carry_f3[2] = {new_rem_carry0[2][55:0], quot_dig0[2][0], 6'b0} = 100100010000000000000000100010000000000000000100000010000000000

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
011111100010101010101010000100010101010101010000101110000000000 + 100100010000000000000000100010000000000000000100000010000000000 = 
000011110010101010101010100110010101010101010100110000000000000
q = 1.001
q ^ 2 = 1.0100010000000000000000000000000000000000000000000000
a_frac - q ^ 2 = 10101001100101010101010101001100101010101010101001100 - 10100010000000000000000000000000000000000000000000000 = 
00000111100101010101010101001100101010101010101001100

// ================================================================================================================================================
// iter[1]:
// ================================================================================================================================================
rem_sum_f3 = 011111100010101010101010000100010101010101010000101110000000000
rem_carry_f3 = 100100010000000000000000100010000000000000000100000010000000000

raw_mask_f3 = 100000000000000000
quot_f3 = 1001000000000000000000000000000000000000000000000000000
quot_m1_f3 = 1000000000000000000000000000000000000000000000000000000

mask_f3[0] = 11110000000000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
11110000000000000000000000000000000000000000000000000000 ^ 
11111000000000000000000000000000000000000000000000000000 = 
00001000000000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0000100000000000000000000000000000000000000000000000000 |
0001000000000000000000000000000000000000000000000000000 = 
0001100000000000000000000000000000000000000000000000000

mask_f3[1] 		= 11111000000000000000000000000000000000000000000000000000
msk_dig[1] 		= 00000100000000000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0000110000000000000000000000000000000000000000000000000

mask_f3[2] 		= 11111100000000000000000000000000000000000000000000000000
msk_dig[2] 		= 00000010000000000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0000011000000000000000000000000000000000000000000000000


rem_sum_f3[62:60] = 011
rem_carry_f3[62:60] = 100
-> 
quot_dig0[0] = 00
->
prev_quot[0] = quot_f3 = 1001000000000000000000000000000000000000000000000000000
prev_quot_m1[0] = quot_m1_f3 = 1000000000000000000000000000000000000000000000000000000
new_quot0_f3[0] = prev_quot[0] & mask_f3[0][55:1] = 1001000000000000000000000000000000000000000000000000000
new_quot0_m1_f3[0] = prev_quot_m1[i] & mask_f3[0][55:1] | msk_dig[0][55:1] = 1000100000000000000000000000000000000000000000000000000

csa_val0[0] = 000000000000000000000000000000000000000000000000000
csa_mux[0] = 000000000000000000000000000000000000000000000000000000000

rem_sum_in[0] = rem_sum_f3[61:0] = 11111100010101010101010000100010101010101010000101110000000000
rem_carry_in[0] = rem_carry_f3[61:0] = 00100010000000000000000100010000000000000000100000010000000000

rem_sum_in[0][61:56] 		= 111111
rem_carry_in[0][61:56] 		= 001000

rem0_sum_zero[0][5:0] 		= 010111
rem0_carry_zero[0][5:0] 	= 110000
rem_sum_msb0[0][5:0] 		= 010111
rem_carry_msb0[0][5:0] 		= 110000

rem_sum_xor[0][56:0] = 
000101010101010100001000101010101010100001011100000000000 ^ 
100000000000000001000100000000000000001000000100000000000 ^ 
000000000000000000000000000000000000000000000000000000000 = 
100101010101010101001100101010101010101001011000000000000
rem_carry_andor[0][57:0] = 0000000000000000000000000000000000000000000001000000000000

new_rem_sum0[0][56:0] = {rem_sum_msb0[0][5:0], rem_sum_xor[0][56: 6]} = 010111100101010101010101001100101010101010101001011000000
new_rem_sum_f3[0] = {new_rem_sum0[0][56:0], 6'b0} = 010111100101010101010101001100101010101010101001011000000000000
new_rem_carry0[0][55:0] = {rem_carry_msb0[0][5:1], rem_carry_andor[0][57: 7]} = 11000000000000000000000000000000000000000000000000100000
new_rem_carry_f3[0] = {new_rem_carry0[0][55:0], quot_dig0[0][0], 6'b0} = 110000000000000000000000000000000000000000000000001000000000000


// ====================================
rem_sum_in[1] = new_rem_sum_f3[0][61:0] = 10111100101010101010101001100101010101010101001011000000000000
rem_carry_in[1] = new_rem_carry_f3[0][61:0] = 10000000000000000000000000000000000000000000000001000000000000

rem_sum_msb0[0][5:3] = 010
rem_carry_msb0[0][5:3] = 110
->
quot_dig0[1] = 01
->
prev_quot[1] = new_quot0_f3[0] = 1001000000000000000000000000000000000000000000000000000
prev_quot_m1[1] = new_quot0_m1_f3[0] = 1000100000000000000000000000000000000000000000000000000
new_quot0_f3[1] = prev_quot[1] & mask_f3[1][55:1] | msk_dig[1][55:1] = 1001010000000000000000000000000000000000000000000000000
new_quot0_m1_f3[1] = prev_quot[1] & mask_f3[1][55:1] = 1001000000000000000000000000000000000000000000000000000

csa_minus_val_sqrt0[1] = {new_quot0_f3[0][53:1], 2'b0} | msk_dig[1][55: 1] = 
0010000000000000000000000000000000000000000000000000000 | 
0000010000000000000000000000000000000000000000000000000 = 
0010010000000000000000000000000000000000000000000000000
csa_val0[1] = ~csa_minus_val0[1][50:0] = 101111111111111111111111111111111111111111111111111
csa_mux[1] = 101111111111111111111111111111111111111111111111111000000

rem_sum_in[1][61:56] 		= 101111
rem_carry_in[1][61:56] 		= 100000
csa_minus_val0[1][54:51] 	=   0010 -> 1101
rem0_sum_minus[1][5:0] 		= 000010
rem0_carry_minus[1][5:0] 	= 111010
rem_sum_msb0[1][5:0] 		= 000010
rem_carry_msb0[1][5:0] 		= 111010

rem_sum_xor[1][56:0] = 
001010101010101010011001010101010101010010110000000000000 ^ 
000000000000000000000000000000000000000000010000000000000 ^ 
101111111111111111111111111111111111111111111111111000000 = 
100101010101010101100110101010101010101101011111111000000
rem_carry_andor[1][57:0] = 0010101010101010100110010101010101010100101100000000000001

new_rem_sum0[1][56:0] = {rem_sum_msb0[1][5:0], rem_sum_xor[1][56: 6]} = 000010100101010101010101100110101010101010101101011111111
new_rem_sum_f3[1] = {new_rem_sum0[1][56:0], 6'b0} = 000010100101010101010101100110101010101010101101011111111000000
new_rem_carry0[1][55:0] = {rem_carry_msb0[1][5:1], rem_carry_andor[1][57: 7]} = 11101001010101010101010011001010101010101010010110000000
new_rem_carry_f3[1] = {new_rem_carry0[1][55:0], quot_dig0[1][0], 6'b0} = 111010010101010101010100110010101010101010100101100000001000000

此时:
new_rem_sum_f3[1] + new_rem_carry_f3[1] = 
000010100101010101010101100110101010101010101101011111111000000 +
111010010101010101010100110010101010101010100101100000001000000 = 
111100111010101010101010011001010101010101010011000000000000000 < 0
q_real = 1.00100
q_real ^ 2 = 1.0100010000000000000000000000000000000000000000000000
a_frac = 1.0101001100101010101010101001100101010101010101001100
diff = 0.0000111100101010101010101001100101010101010101001100

{new_quot0_m1_f3[1], 1'b0} | msk_dig[2] = 
10010000000000000000000000000000000000000000000000000000 |
00000010000000000000000000000000000000000000000000000000 =
10010010000000000000000000000000000000000000000000000000
{1'b0, ({new_quot0_m1_f3[1], 1'b0} | msk_dig[2]), 6'b0} = 010010010000000000000000000000000000000000000000000000000000000
111100111010101010101010011001010101010101010011000000000000000 +
010010010000000000000000000000000000000000000000000000000000000 = 
001111001010101010101010011001010101010101010011000000000000000
00000111100101010101010101001100101010101010101001100

// ====================================
rem_sum_in[2] = new_rem_sum_f3[1][61:0] = 00010100101010101010101100110101010101010101101011111111000000
rem_carry_in[2] = new_rem_carry_f3[1][61:0] = 11010010101010101010100110010101010101010100101100000001000000

rem_sum_msb0[1][5:3] = 000
rem_carry_msb0[1][5:3] = 111
->
quot_dig0[2] = 00
->
prev_quot[2] = new_quot0_f3[1] = 1001010000000000000000000000000000000000000000000000000
prev_quot_m1[2] = new_quot0_m1_f3[1] = 1001000000000000000000000000000000000000000000000000000
new_quot0_f3[2] = prev_quot[2] & mask_f3[2][55:1] = 1001010000000000000000000000000000000000000000000000000
new_quot0_m1_f3[2] = prev_quot_m1[2] & mask_f3[2][55:1] | msk_dig[2][55:1] = 1001001000000000000000000000000000000000000000000000000

csa_val0[2] = csa_plus_val0[2][50:0] = 000000000000000000000000000000000000000000000000000
csa_mux[1] = 000000000000000000000000000000000000000000000000000000000

rem_sum_in[2][61:56] 		= 000101
rem_carry_in[2][61:56] 		= 110100

rem0_sum_zero[2][5:0] 		= 010001
rem0_carry_zero[2][5:0] 	= 101000
rem_sum_msb0[2][5:0] 		= 010001
rem_carry_msb0[2][5:0] 		= 101000

rem_sum_xor[2][56:0] = 
001010101010101011001101010101010101011010111111110000000 ^ 
101010101010101001100101010101010101001011000000010000000 ^ 
000000000000000000000000000000000000000000000000000000000 = 
100000000000000010101000000000000000010001111111100000000
rem_carry_andor[2][57:0] = 0010101010101010010001010101010101010010100000000100000000

new_rem_sum0[2][56:0] = {rem_sum_msb0[2][5:0], rem_sum_xor[2][56: 6]} = 010001100000000000000010101000000000000000010001111111100
new_rem_sum_f3[2] = {new_rem_sum0[2][56:0], 6'b0} = 010001100000000000000010101000000000000000010001111111100000000
new_rem_carry0[2][55:0] = {rem_carry_msb0[2][5:1], rem_carry_andor[2][57: 7]} = 10100001010101010101001000101010101010101001010000000010
new_rem_carry_f3[2] = {new_rem_carry0[2][55:0], quot_dig0[2][0], 6'b0} = 101000010101010101010010001010101010101010010100000000100000000

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
010001100000000000000010101000000000000000010001111111100000000 +
101000010101010101010010001010101010101010010100000000100000000 = 
111001110101010101010100110010101010101010100110000000000000000 < 0
q_real = 1.001_001
q_real ^ 2 = 1.0100110100010000000000000000000000000000000000000000
a_frac - q ^ 2 = 10101001100101010101010101001100101010101010101001100 - 10100110100010000000000000000000000000000000000000000 = 
0.0000011000011010101010101001100101010101010101001100

// 下个iter中: 
msk_dig[0] = 00000001000000000000000000000000000000000000000000000000
{new_quot0_m1_f3[2], 1'b0} | msk_dig[0] = 
10010010000000000000000000000000000000000000000000000000 |
00000001000000000000000000000000000000000000000000000000 = 
10010011000000000000000000000000000000000000000000000000
{1'b0, ({new_quot0_m1_f3[2], 1'b0} | msk_dig[0]), 6'b0} = 
010010011000000000000000000000000000000000000000000000000000000

111001110101010101010100110010101010101010100110000000000000000 + 
010010011000000000000000000000000000000000000000000000000000000 = 
001100001101010101010100110010101010101010100110000000000000000





// ================================================================================================================================================
对fp16[15:0].sqrt来一个.....
a_frac = 1.1010001100
sqrt(a_frac << 1) = 1.1100111100_1_0101111110...
init_rem_sum_adj[14:0] = 010010001100000
// ================================================================================================================================================
// iter[0]:
// ================================================================================================================================================
rem_sum_f3[14:0] = 010010001100000
rem_carry_f3[14:0] = 000000000000000

quot_f3[12:0] = 1000000000000
quot_m1_f3[12:0] = 0000000000000

raw_mask_f3 = 000000000000000000
mask_f3[0] = 10000000000000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
10000000000000000000000000000000000000000000000000000000 ^ 
11000000000000000000000000000000000000000000000000000000 = 
01000000000000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0100000000000000000000000000000000000000000000000000000 |
1000000000000000000000000000000000000000000000000000000 = 
1100000000000000000000000000000000000000000000000000000

mask_f3[1] 		= 11000000000000000000000000000000000000000000000000000000
msk_dig[1] 		= 00100000000000000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0110000000000000000000000000000000000000000000000000000

mask_f3[2] 		= 11100000000000000000000000000000000000000000000000000000
msk_dig[2] 		= 00010000000000000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0011000000000000000000000000000000000000000000000000000

rem_sum_f3[14:12] = 010
rem_carry_f3[14:12] = 000
-> 
quot_dig3[0] = 01
->
prev_quot[0][12:0] = quot_f3[12:0] = 1000000000000
prev_quot_m1[0] = quot_m1_f3[12:0] = 0000000000000
new_quot3_f3[0] = prev_quot[0] & mask_f3[0][55:43] | msk_dig[0][55:43] = 1100000000000
new_quot3_m1_f3[0] = prev_quot[0] & mask_f3[0][55:43] = 1000000000000

csa_minus_val_sqrt3[0] = {quot_f3[11: 1], 1'b0} | msk_dig[0][55:44] = 
000000000000 | 
010000000000 = 
010000000000
csa_minus_val3[0] = {2'b00, csa_minus_val_sqrt3[0]} = 00010000000000
csa_val3[0] = ~csa_minus_val3[0][13:0] = 11101111111111
csa_mux[0][14:0] = {csa_val3[0][13:0], 1'b0} = 111011111111110

rem_sum_in[0][13:0] = rem_sum_f3[13:0] = 10010001100000
rem_carry_in[0][13:0] = rem_carry_f3[13:0] = 00000000000000

rem_sum_in[0][13:8] 		= 100100
rem_carry_in[0][13:8] 		= 000000
csa_minus_val3[0][11:8] 	=   0100 -> 1011
rem3_sum_minus[0][5:0] 		= 001111
rem3_carry_minus[0][5:0] 	= 000001
rem_sum_msb3[0][5:0] 		= 001111
rem_carry_msb3[0][5:0] 		= 000001

rem_sum_xor[0][9:0] = 
0011000000 ^ 
0000000000 ^ 
1111111110 = 
1100111110
rem_carry_andor[0][10:0] = 00110000001

new_rem_sum3[0][13:0] = {rem_sum_msb3[0][5:0], rem_sum_xor[0][ 8: 1]} = 00111110011111
new_rem_sum_f3[0] = {new_rem_sum3[0][13: 0], 1'b0} = 001111100111110
new_rem_carry3[0][12:0] = {rem_carry_msb3[0][5:1], rem_carry_andor[0][ 9: 2]} = 0000001100000
new_rem_carry_f3[0] = {new_rem_carry3[0][12: 0], quot_dig3[0][0], 1'b0} = 000000110000010


此时:
new_rem_sum_f3[0] + new_rem_carry_f3[0] = 
001111100111110 + 
000000110000010 = 
010000011000000

q_real = 1.1
q_real ^ 2 = 10.01
a_frac << 1 = 11.0100011000
diff = 1.0000011000000000

// ======================
rem_sum_in[1] = new_rem_sum_f3[0][14:0] = 001111100111110
rem_carry_in[1] = new_rem_carry_f3[0][14:0] = 000000110000010

rem_sum_msb3[0][5:3] = 001
rem_carry_msb3[0][5:3] = 000
->
quot_dig3[1] = 01
->
prev_quot[1] = new_quot3_f3[0] = 1100000000000
prev_quot_m1[1] = new_quot3_m1_f3[0] = 1000000000000
new_quot3_f3[1] = prev_quot[1] & mask_f3[1][55:43] | msk_dig[1][55:43] = 1110000000000
new_quot3_m1_f3[1] = prev_quot[1] & mask_f3[1][55:43] = 1100000000000

csa_minus_val_sqrt3[1] = {new_quot3_f3[0][11: 1], 1'b0} | msk_dig[1][55:44] = 
100000000000 | 
001000000000 = 
101000000000
csa_minus_val3[1] = {2'b00, csa_minus_val_sqrt3[1]} = 00101000000000
csa_val3[1] = ~csa_minus_val3[1][13:0] = 11010111111111
csa_mux[1][14:0] = {csa_val3[1][13:0], 1'b0} = 110101111111110

rem_sum_in[1][13:0] = 01111100111110
rem_carry_in[1][13:0] = 00000110000010

rem_sum_in[1][13:8] 		= 011111
rem_carry_in[1][13:8] 		= 000001
csa_minus_val3[1][11:8] 	=   1010 -> 0101
rem3_sum_minus[1][5:0] 		= 011011
rem3_carry_minus[1][5:0] 	= 101011
rem_sum_msb3[1][5:0] 		= 011011
rem_carry_msb3[1][5:0] 		= 101011

rem_sum_xor[1][9:0] = 
1001111100 ^ 
1100000100 ^ 
1111111110 = 
1010000110
rem_carry_andor[1][10:0] = 11011111001

new_rem_sum3[1][13:0] = {rem_sum_msb3[1][5:0], rem_sum_xor[1][ 8: 1]} = 01101101000011
new_rem_sum_f3[1] = {new_rem_sum3[1][13: 0], 1'b0} = 011011010000110
new_rem_carry3[1][12:0] = {rem_carry_msb3[1][5:1], rem_carry_andor[1][ 9: 2]} = 1010110111110
new_rem_carry_f3[1] = {new_rem_carry3[1][12: 0], quot_dig3[1][0], 1'b0} = 101011011111010

此时:
new_rem_sum_f3[1] + new_rem_carry_f3[1] = 
011011010000110 + 
101011011111010 = 
000110110000000

q_real = 1.11
q_real ^ 2 = 11.00010000
a_frac << 1 = 11.0100011000
diff = 0.001101100000000

// ======================
rem_sum_in[2] = new_rem_sum_f3[1][14:0] = 011011010000110
rem_carry_in[2] = new_rem_carry_f3[1][14:0] = 101011011111010

rem_sum_msb3[1][5:3] = 011
rem_carry_msb3[1][5:3] = 101
->
quot_dig3[2] = 01
->
prev_quot[2] = new_quot3_f3[1] = 1110000000000
prev_quot_m1[2] = new_quot3_m1_f3[1] = 1100000000000
new_quot3_f3[2] = prev_quot[2] & mask_f3[2][55:43] | msk_dig[2][55:43] = 1111000000000
new_quot3_m1_f3[2] = prev_quot[2] & mask_f3[2][55:43] = 1110000000000

csa_minus_val_sqrt3[2] = {new_quot3_f3[1][11: 1], 1'b0} | msk_dig[2][55:44] = 
110000000000 | 
000100000000 = 
110100000000
csa_minus_val3[2] = {2'b00, csa_minus_val_sqrt3[2]} = 00110100000000
csa_val3[2] = ~csa_minus_val3[2][13:0] = 11001011111111
csa_mux[2][14:0] = {csa_val3[2][13:0], 1'b0} = 110010111111110

rem_sum_in[2][13:0] = 11011010000110
rem_carry_in[2][13:0] = 01011011111010

rem_sum_in[2][13:8] 		= 110110
rem_carry_in[2][13:8] 		= 010110
csa_minus_val3[2][11:8] 	=   1101 -> 0010
rem3_sum_minus[2][5:0] 		= 000010
rem3_carry_minus[2][5:0] 	= 101101
rem_sum_msb3[2][5:0] 		= 000010
rem_carry_msb3[2][5:0] 		= 101101

rem_sum_xor[2][9:0] = 
0100001100 ^ 
0111110100 ^ 
0111111110 = 
0100000110
rem_carry_andor[2][10:0] = 01111111001
new_rem_sum3[2][13:0] = {rem_sum_msb3[2][5:0], rem_sum_xor[2][ 8: 1]} = 00001010000011
new_rem_sum_f3[2] = {new_rem_sum3[2][13: 0], 1'b0} = 000010100000110
new_rem_carry3[2][12:0] = {rem_carry_msb3[2][5:1], rem_carry_andor[2][ 9: 2]} = 1011011111110
new_rem_carry_f3[2] = {new_rem_carry3[2][12: 0], quot_dig3[2][0], 1'b0} = 101101111111010

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
000010100000110 + 
101101111111010 = 
110000100000000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
下次迭代: msk_dig[0][55:42] = 00001000000000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[2], 1'b0} | 00001000000000} = 011101000000000
110000100000000 + 
011101000000000 = 
001101100000000

q_real = 1.110
q_real ^ 2 = 11.00010000
a_frac << 1 = 11.0100011000
diff = 0.0011011000000000

// ================================================================================================================================================
// iter[1]:
// ================================================================================================================================================
rem_sum_f3[14:0] = 000010100000110
rem_carry_f3[14:0] = 101101111111010

quot_f3[12:0] = 1111000000000
quot_m1_f3[12:0] = 1110000000000

raw_mask_f3 = 100000000000000000
mask_f3[0] = 11110000000000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
11110000000000000000000000000000000000000000000000000000 ^ 
11111000000000000000000000000000000000000000000000000000 = 
00001000000000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0000100000000000000000000000000000000000000000000000000 |
0001000000000000000000000000000000000000000000000000000 = 
0001100000000000000000000000000000000000000000000000000

mask_f3[1] 		= 11111000000000000000000000000000000000000000000000000000
msk_dig[1] 		= 00000100000000000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0000110000000000000000000000000000000000000000000000000

mask_f3[2] 		= 11111100000000000000000000000000000000000000000000000000
msk_dig[2] 		= 00000010000000000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0000011000000000000000000000000000000000000000000000000

rem_sum_f3[14:12] = 000
rem_carry_f3[14:12] = 101
-> 
quot_dig3[0] = 10
->
prev_quot[0][12:0] = quot_f3[12:0] = 1111000000000
prev_quot_m1[0] = quot_m1_f3[12:0] = 1110000000000
new_quot3_f3[0] = prev_quot_m1[0] & mask_f3[0][55:43] | msk_dig[0][55:43] = 1110100000000
new_quot3_m1_f3[0] = prev_quot_m1[0] & mask_f3[0][55:43] = 1110000000000

csa_plus_val_sqrt3[0] = {quot_m1_f3[11: 1], 1'b0} | msk_dig_3[0][54:43] = 
110000000000 | 
000110000000 = 
110110000000
csa_plus_val3[0] = {2'b00, csa_plus_val_sqrt3[0]} = 00110110000000
csa_val3[0] = csa_plus_val3[0][13:0] = 00110110000000
csa_mux[0][14:0] = {csa_val3[0][13:0], 1'b0} = 001101100000000

rem_sum_in[0][13:0] = rem_sum_f3[13:0] = 00010100000110
rem_carry_in[0][13:0] = rem_carry_f3[13:0] = 01101111111010

rem_sum_in[0][13:8] 		= 000101
rem_carry_in[0][13:8] 		= 011011
csa_plus_val3[0][11:8] 		=   1101
rem3_sum_plus[0][5:0] 		= 000011
rem3_carry_plus[0][5:0] 	= 111010
rem_sum_msb3[0][5:0] 		= 000011
rem_carry_msb3[0][5:0] 		= 111010

rem_sum_xor[0][9:0] = 
1000001100 ^ 
1111110100 ^ 
1100000000 = 
1011111000
rem_carry_andor[0][10:0] = 11000001001

new_rem_sum3[0][13:0] = {rem_sum_msb3[0][5:0], rem_sum_xor[0][ 8: 1]} = 00001101111100
new_rem_sum_f3[0] = {new_rem_sum3[0][13: 0], 1'b0} = 000011011111000
new_rem_carry3[0][12:0] = {rem_carry_msb3[0][5:1], rem_carry_andor[0][ 9: 2]} = 1110110000010
new_rem_carry_f3[0] = {new_rem_carry3[0][12: 0], quot_dig3[0][0], 1'b0} = 111011000001000


此时:
new_rem_sum_f3[0] + new_rem_carry_f3[0] = 
000011011111000 + 
111011000001000 = 
111110100000000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[1][55:42] = 00000100000000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[0], 1'b0} | 00000100000000} = 011100100000000
111110100000000 + 
011100100000000 = 
011011000000000

q_real = 1.1100
q_real ^ 2 = 11.00010000
a_frac << 1 = 11.0100011000
diff = 0.0011011000000000

// ======================
rem_sum_in[1] = new_rem_sum_f3[0][14:0] = 000011011111000
rem_carry_in[1] = new_rem_carry_f3[0][14:0] = 111011000001000

rem_sum_msb3[0][5:3] = 000
rem_carry_msb3[0][5:3] = 111
->
quot_dig3[1] = 00
->
prev_quot[1] = new_quot3_f3[0] = 1110100000000
prev_quot_m1[1] = new_quot3_m1_f3[0] = 1110000000000
new_quot3_f3[1] = prev_quot[1] & mask_f3[1][55:43] = 1110100000000
new_quot3_m1_f3[1] = prev_quot_m1[1] & mask_f3[1][55:43] | msk_dig[1][55:43] = 1110010000000

// Not used...
// csa_minus_val_sqrt3[1] = {new_quot3_f3[0][11: 1], 1'b0} | msk_dig[1][55:44] = 
// 100000000000 | 
// 001000000000 = 
// 101000000000
// csa_minus_val3[1] = {2'b00, csa_minus_val_sqrt3[1]} = 00101000000000
csa_val3[1] = 00000000000000
csa_mux[1][14:0] = {csa_val3[1][13:0], 1'b0} = 000000000000000

rem_sum_in[1][13:0] = 00011011111000
rem_carry_in[1][13:0] = 11011000001000

rem_sum_in[1][13:8] 		= 000110
rem_carry_in[1][13:8] 		= 110110
// csa_minus_val3[1][11:8] 	=   1010 -> 0101
rem3_sum_zero[1][5:0] 		= 010000
rem3_carry_zero[1][5:0] 	= 101100
rem_sum_msb3[1][5:0] 		= 010000
rem_carry_msb3[1][5:0] 		= 101100


rem_sum_xor[1][9:0] = 
0111110000 ^ 
0000010000 ^ 
0000000000 = 
0111100000
rem_carry_andor[1][10:0] = 00000100000

new_rem_sum3[1][13:0] = {rem_sum_msb3[1][5:0], rem_sum_xor[1][ 8: 1]} = 01000011110000
new_rem_sum_f3[1] = {new_rem_sum3[1][13: 0], 1'b0} = 010000111100000
new_rem_carry3[1][12:0] = {rem_carry_msb3[1][5:1], rem_carry_andor[1][ 9: 2]} = 1011000001000
new_rem_carry_f3[1] = {new_rem_carry3[1][12: 0], quot_dig3[1][0], 1'b0} = 101100000100000

此时:
new_rem_sum_f3[1] + new_rem_carry_f3[1] = 
010000111100000 + 
101100000100000 = 
111101000000000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[2][55:42] = 00000010000000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[1], 1'b0} | 00000010000000} = 011100110000000
111101000000000 + 
011100110000000 = 
011001110000000

q_real = 1.11001
q_real ^ 2 = 11.001011000100
a_frac << 1 = 11.0100011000
diff = 0.0001100111000000

// ======================
rem_sum_in[2] = new_rem_sum_f3[1][14:0] = 010000111100000
rem_carry_in[2] = new_rem_carry_f3[1][14:0] = 101100000100000

rem_sum_msb3[1][5:3] = 010
rem_carry_msb3[1][5:3] = 101
->
quot_dig3[2] = 00
->
prev_quot[2] = new_quot3_f3[1] = 1110100000000
prev_quot_m1[2] = new_quot3_m1_f3[1] = 1110010000000
new_quot3_f3[2] = prev_quot[2] & mask_f3[2][55:43] = 1110100000000
new_quot3_m1_f3[2] = prev_quot_m1[2] & mask_f3[2][55:43] | msk_dig[2][55:43] = 1110011000000

// Not used...
// csa_minus_val_sqrt3[2] = {new_quot3_f3[1][11: 1], 1'b0} | msk_dig[2][55:44] = 
// 110000000000 | 
// 000100000000 = 
// 110100000000
// csa_minus_val3[2] = {2'b00, csa_minus_val_sqrt3[2]} = 00110100000000
csa_val3[2] = 0000000000000
csa_mux[2][14:0] = {csa_val3[2][13:0], 1'b0} = 00000000000000

rem_sum_in[2][13:0] = 10000111100000
rem_carry_in[2][13:0] = 01100000100000

rem_sum_in[2][13:8] 		= 100001
rem_carry_in[2][13:8] 		= 011000
// csa_minus_val3[2][11:8] 	=   1101 -> 0010
rem3_sum_zero[2][5:0] 		= 011001
rem3_carry_zero[2][5:0] 	= 100000
rem_sum_msb3[2][5:0] 		= 011001
rem_carry_msb3[2][5:0] 		= 100000

rem_sum_xor[2][9:0] = 
1111000000 ^ 
0001000000 ^ 
0000000000 = 
1110000000
rem_carry_andor[2][10:0] = 00010000000

new_rem_sum3[2][13:0] = {rem_sum_msb3[2][5:0], rem_sum_xor[2][ 8: 1]} = 01100111000000
new_rem_sum_f3[2] = {new_rem_sum3[2][13: 0], 1'b0} = 011001110000000
new_rem_carry3[2][12:0] = {rem_carry_msb3[2][5:1], rem_carry_andor[2][ 9: 2]} = 1000000100000
new_rem_carry_f3[2] = {new_rem_carry3[2][12: 0], quot_dig3[2][0], 1'b0} = 100000010000000

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
011001110000000 + 
100000010000000 = 
111010000000000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
下次迭代: msk_dig[0][55:42] = 00000001000000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[2], 1'b0} | 00000001000000} = 011100111000000
111010000000000 + 
011100111000000 = 
010110111000000

q_real = 1.110011
q_real ^ 2 = 11.001110101001000
a_frac << 1 = 11.0100011000
diff = 0.000010110111000

// ================================================================================================================================================
// iter[2]:
// ================================================================================================================================================
rem_sum_f3[14:0] = 011001110000000
rem_carry_f3[14:0] = 100000010000000

quot_f3[12:0] = 1110100000000
quot_m1_f3[12:0] = 1110011000000

raw_mask_f3 = 11000000000000000
mask_f3[0] = 11111110000000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
11111110000000000000000000000000000000000000000000000000 ^ 
11111111000000000000000000000000000000000000000000000000 = 
00000001000000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0000000100000000000000000000000000000000000000000000000 |
0000001000000000000000000000000000000000000000000000000 = 
0000001100000000000000000000000000000000000000000000000

mask_f3[1] 		= 11111111000000000000000000000000000000000000000000000000
msk_dig[1] 		= 00000000100000000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0000000110000000000000000000000000000000000000000000000

mask_f3[2] 		= 11111111100000000000000000000000000000000000000000000000
msk_dig[2] 		= 00000000010000000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0000000011000000000000000000000000000000000000000000000

rem_sum_f3[14:12] = 011
rem_carry_f3[14:12] = 100
-> 
quot_dig3[0] = 00
->
prev_quot[0][12:0] = quot_f3[12:0] = 1110100000000
prev_quot_m1[0] = quot_m1_f3[12:0] = 1110011000000
new_quot3_f3[0] = prev_quot[0] & mask_f3[0][55:43] = 1110100000000
new_quot3_m1_f3[0] = prev_quot_m1[0] & mask_f3[0][55:43] | msk_dig[0][55:43] = 1110011100000

// Not used...
// csa_plus_val_sqrt3[0] = {quot_m1_f3[11: 1], 1'b0} | msk_dig_3[0][54:43] = 
// 110000000000 | 
// 0001100000000 = 
// 110110000000
// csa_plus_val3[0] = {2'b00, csa_plus_val_sqrt3[0]} = 00110110000000
csa_val3[0] = 00000000000000
csa_mux[0][14:0] = {csa_val3[0][13:0], 1'b0} = 000000000000000

rem_sum_in[0][13:0] = rem_sum_f3[13:0] = 11001110000000
rem_carry_in[0][13:0] = rem_carry_f3[13:0] = 00000010000000

rem_sum_in[0][13:8] 		= 110011
rem_carry_in[0][13:8] 		= 000000
// csa_plus_val3[0][11:8] 		=   1101
rem3_sum_zero[0][5:0] 		= 010011
rem3_carry_zero[0][5:0] 	= 100000
rem_sum_msb3[0][5:0] 		= 010011
rem_carry_msb3[0][5:0] 		= 100000

rem_sum_xor[0][9:0] = 
1100000000 ^ 
0100000000 ^ 
0000000000 = 
1000000000
rem_carry_andor[0][10:0] = 01000000000

new_rem_sum3[0][13:0] = {rem_sum_msb3[0][5:0], rem_sum_xor[0][ 8: 1]} = 01001100000000
new_rem_sum_f3[0] = {new_rem_sum3[0][13: 0], 1'b0} = 010011000000000
new_rem_carry3[0][12:0] = {rem_carry_msb3[0][5:1], rem_carry_andor[0][ 9: 2]} = 1000010000000
new_rem_carry_f3[0] = {new_rem_carry3[0][12: 0], quot_dig3[0][0], 1'b0} = 100001000000000


此时:
new_rem_sum_f3[0] + new_rem_carry_f3[0] = 
010011000000000 + 
100001000000000 = 
110100000000000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[1][55:42] = 00000000100000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[0], 1'b0} | 00000000100000} = 011100111100000
110100000000000 + 
011100111100000 = 
010000111100000

q_real = 1.1100111
q_real ^ 2 = 11.00010000
a_frac << 1 = 11.0100011000
diff = 0.00000100001111000000

// ======================
rem_sum_in[1] = new_rem_sum_f3[0][14:0] = 010011000000000
rem_carry_in[1] = new_rem_carry_f3[0][14:0] = 100001000000000

rem_sum_msb3[0][5:3] = 010
rem_carry_msb3[0][5:3] = 100
->
quot_dig3[1] = 10
->
prev_quot[1] = new_quot3_f3[0] = 1110100000000
prev_quot_m1[1] = new_quot3_m1_f3[0] = 1110011100000
new_quot3_f3[1] = prev_quot_m1[1] & mask_f3[1][55:43] | msk_dig[1][55:43] = 1110011110000
new_quot3_m1_f3[1] = prev_quot_m1[1] & mask_f3[1][55:43] = 1110011100000

csa_plus_val_sqrt3[1] = {new_quot3_m1_f3[0][11:1], 1'b0} | msk_dig_3[1][54:43] = 
110011100000 | 
000000011000 = 
110011111000
csa_plus_val3[1] = {2'b00, csa_plus_val_sqrt3[1]} = 00110011111000
csa_val3[1] = csa_plus_val3[1][13:0] = 00110011111000
csa_mux[1][14:0] = {csa_val3[1][13:0], 1'b0} = 001100111110000


rem_sum_in[1][13:0] = 10011000000000
rem_carry_in[1][13:0] = 00001000000000

rem_sum_in[1][13:8] 		= 100110
rem_carry_in[1][13:8] 		= 000010
csa_plus_val3[1][11:8] 		=   1100
rem3_sum_plus[1][5:0] 		= 011000
rem3_carry_plus[1][5:0] 	= 101100
rem_sum_msb3[1][5:0] 		= 011000
rem_carry_msb3[1][5:0] 		= 101100

rem_sum_xor[1][9:0] = 
0000000000 ^ 
0000000000 ^ 
0111110000 = 
0111110000
rem_carry_andor[1][10:0] = 00000000000

new_rem_sum3[1][13:0] = {rem_sum_msb3[1][5:0], rem_sum_xor[1][ 8: 1]} = 01100011111000
new_rem_sum_f3[1] = {new_rem_sum3[1][13: 0], 1'b0} = 011000111110000
new_rem_carry3[1][12:0] = {rem_carry_msb3[1][5:1], rem_carry_andor[1][ 9: 2]} = 1011000000000
new_rem_carry_f3[1] = {new_rem_carry3[1][12: 0], quot_dig3[1][0], 1'b0} = 101100000000000

此时:
new_rem_sum_f3[1] + new_rem_carry_f3[1] = 
011000111110000 + 
101100000000000 = 
000100111110000

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[2][55:42] = 00000000010000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[1], 1'b0} | 00000000010000} = 011100111010000
// 111101000000000 + 
// 011100110000000 = 
// 011001110000000

q_real = 1.11001111
q_real ^ 2 = 11.01000101011000010
a_frac << 1 = 11.0100011000
diff = 0.0000000010011111000000

// ======================
rem_sum_in[2] = new_rem_sum_f3[1][14:0] = 011000111110000
rem_carry_in[2] = new_rem_carry_f3[1][14:0] = 101100000000000

rem_sum_msb3[1][5:3] = 011
rem_carry_msb3[1][5:3] = 101
->
quot_dig3[2] = 01
->
prev_quot[2] = new_quot3_f3[1] = 1110011110000
prev_quot_m1[2] = new_quot3_m1_f3[1] = 1110011100000
new_quot3_f3[2] = prev_quot[2] & mask_f3[2][55:43] | msk_dig[2][55:43] = 1110011111000
new_quot3_m1_f3[2] = prev_quot[2] & mask_f3[2][55:43] = 1110011110000

csa_minus_val_sqrt3[2] = {new_quot3_f3[1][11: 1], 1'b0} | msk_dig[2][55:44] = 
110011110000 | 
000000000100 = 
110011110100
csa_minus_val3[2] = {2'b00, csa_minus_val_sqrt3[2]} = 00110011110100
csa_val3[2] = ~csa_minus_val3[2][13:0] = 11001100001011
csa_mux[2][14:0] = {csa_val3[2][13:0], 1'b0} = 110011000010110

rem_sum_in[2][13:0] = 11000111110000
rem_carry_in[2][13:0] = 01100000000000

rem_sum_in[2][13:8] 		= 110001
rem_carry_in[2][13:8] 		= 011000
csa_minus_val3[2][11:8] 	=   1100 -> 0011
rem3_sum_minus[2][5:0] 		= 001010
rem3_carry_minus[2][5:0] 	= 100011
rem_sum_msb3[2][5:0] 		= 001010
rem_carry_msb3[2][5:0] 		= 100011

rem_sum_xor[2][9:0] = 
1111100000 ^ 
0000000000 ^ 
1000010110 = 
0111110110
rem_carry_andor[2][10:0] = 10000000001

new_rem_sum3[2][13:0] = {rem_sum_msb3[2][5:0], rem_sum_xor[2][ 8: 1]} = 00101011111011
new_rem_sum_f3[2] = {new_rem_sum3[2][13: 0], 1'b0} = 001010111110110
new_rem_carry3[2][12:0] = {rem_carry_msb3[2][5:1], rem_carry_andor[2][ 9: 2]} = 1000100000000
new_rem_carry_f3[2] = {new_rem_carry3[2][12: 0], quot_dig3[2][0], 1'b0} = 100010000000010

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
001010111110110 + 
100010000000010 = 
101100111111000


// TODO: 恢复余数的方法只是自己根据fp64猜的...
下次迭代: msk_dig[0][55:42] = 00000000001000
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[2], 1'b0} | 00000000001000} = 011100111101000
101100111111000 + 
011100111101000 = 
001001111100000

q_real = 1.110011110
q_real ^ 2 = 11.01000101011000010
a_frac << 1 = 11.0100011000
diff = 0.000000001001111100000


// ================================================================================================================================================
// iter[3]:
// ================================================================================================================================================
rem_sum_f3[14:0] = 001010111110110
rem_carry_f3[14:0] = 100010000000010

quot_f3[12:0] = 1110011111000
quot_m1_f3[12:0] = 1110011110000

raw_mask_f3 = 11100000000000000
mask_f3[0] = 11111111110000000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
11111111110000000000000000000000000000000000000000000000 ^ 
11111111111000000000000000000000000000000000000000000000 = 
00000000001000000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0000000000100000000000000000000000000000000000000000000 |
0000000001000000000000000000000000000000000000000000000 = 
0000000001100000000000000000000000000000000000000000000

mask_f3[1] 		= 11111111111000000000000000000000000000000000000000000000
msk_dig[1] 		= 00000000000100000000000000000000000000000000000000000000
msk_dig_3[1] 	= 0000000000110000000000000000000000000000000000000000000

mask_f3[2] 		= 11111111111100000000000000000000000000000000000000000000
msk_dig[2] 		= 00000000000010000000000000000000000000000000000000000000
msk_dig_3[2] 	= 0000000000011000000000000000000000000000000000000000000

rem_sum_f3[14:12] = 001
rem_carry_f3[14:12] = 100
-> 
quot_dig3[0] = 10
->
prev_quot[0][12:0] = quot_f3[12:0] = 1110011111000
prev_quot_m1[0] = quot_m1_f3[12:0] = 1110011110000
new_quot3_f3[0] = prev_quot_m1[0] & mask_f3[0][55:43] | msk_dig[0][55:43] = 1110011110100
new_quot3_m1_f3[0] = prev_quot_m1[0] & mask_f3[0][55:43] = 1110011110000

csa_plus_val_sqrt3[0] = {quot_m1_f3[11: 1], 1'b0} | msk_dig_3[0][54:43] = 
110011110000 | 
000000000110 = 
110011110110
csa_plus_val3[0] = {2'b00, csa_plus_val_sqrt3[0]} = 00110011110110
csa_val3[0] = csa_plus_val3[0][13:0] = 00110011110110
csa_mux[0][14:0] = {csa_val3[0][13:0], 1'b0} = 001100111101100

rem_sum_in[0][13:0] = rem_sum_f3[13:0] = 01010111110110
rem_carry_in[0][13:0] = rem_carry_f3[13:0] = 00010000000010

rem_sum_in[0][13:8] 		= 010101
rem_carry_in[0][13:8] 		= 000100
csa_plus_val3[0][11:8] 		=   1100
rem3_sum_plus[0][5:0] 		= 001101
rem3_carry_plus[0][5:0] 	= 101000
rem_sum_msb3[0][5:0] 		= 001101
rem_carry_msb3[0][5:0] 		= 101000

rem_sum_xor[0][9:0] = 
1111101100 ^ 
0000000100 ^ 
0111101100 = 
1000000100
rem_carry_andor[0][10:0] = 01111011000

new_rem_sum3[0][13:0] = {rem_sum_msb3[0][5:0], rem_sum_xor[0][ 8: 1]} = 00110100000010
new_rem_sum_f3[0] = {new_rem_sum3[0][13: 0], 1'b0} = 001101000000100
new_rem_carry3[0][12:0] = {rem_carry_msb3[0][5:1], rem_carry_andor[0][ 9: 2]} = 1010011110110
new_rem_carry_f3[0] = {new_rem_carry3[0][12: 0], quot_dig3[0][0], 1'b0} = 101001111011000


此时:
new_rem_sum_f3[0] + new_rem_carry_f3[0] = 
001101000000100 + 
101001111011000 = 
110110111011100

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[1][55:42] = 00000000000100
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[0], 1'b0} | 00000000000100} = 011100111100100
110110111011100 + 
011100111100100 = 
010011111000000

q_real = 1.1100111100
q_real ^ 2 = 11.0100010101100001000
a_frac << 1 = 11.0100011000
diff = 0.0000000010011111000000

// ======================
rem_sum_in[1] = new_rem_sum_f3[0][14:0] = 001101000000100
rem_carry_in[1] = new_rem_carry_f3[0][14:0] = 101001111011000

rem_sum_msb3[0][5:3] = 001
rem_carry_msb3[0][5:3] = 101
->
quot_dig3[1] = 10
->
prev_quot[1] = new_quot3_f3[0] = 1110011111000
prev_quot_m1[1] = new_quot3_m1_f3[0] = 1110011110000
new_quot3_f3[1] = prev_quot_m1[1] & mask_f3[1][55:43] | msk_dig[1][55:43] = 1110011110010
new_quot3_m1_f3[1] = prev_quot_m1[1] & mask_f3[1][55:43] = 1110011110000

csa_plus_val_sqrt3[1] = {new_quot3_m1_f3[0][11:1], 1'b0} | msk_dig_3[1][54:43] = 
110011110000 | 
000000000011 = 
110011110011
csa_plus_val3[1] = {2'b00, csa_plus_val_sqrt3[1]} = 00110011110011
csa_val3[1] = csa_plus_val3[1][13:0] = 00110011110011
csa_mux[1][14:0] = {csa_val3[1][13:0], 1'b0} = 001100111100110


rem_sum_in[1][13:0] = 01101000000100
rem_carry_in[1][13:0] = 01001111011000

rem_sum_in[1][13:8] 		= 011010
rem_carry_in[1][13:8] 		= 010011
csa_plus_val3[1][11:8] 		=   1100
rem3_sum_plus[1][5:0] 		= 010101
rem3_carry_plus[1][5:0] 	= 110100
rem_sum_msb3[1][5:0] 		= 010101
rem_carry_msb3[1][5:0] 		= 110100

rem_sum_xor[1][9:0] = 
0000001000 ^ 
1110110000 ^ 
0111100110 = 
1001011110
rem_carry_andor[1][10:0] = 01101000000

new_rem_sum3[1][13:0] = {rem_sum_msb3[1][5:0], rem_sum_xor[1][ 8: 1]} = 01010100101111
new_rem_sum_f3[1] = {new_rem_sum3[1][13: 0], 1'b0} = 010101001011110
new_rem_carry3[1][12:0] = {rem_carry_msb3[1][5:1], rem_carry_andor[1][ 9: 2]} = 1101011010000
new_rem_carry_f3[1] = {new_rem_carry3[1][12: 0], quot_dig3[1][0], 1'b0} = 110101101000000

此时:
new_rem_sum_f3[1] + new_rem_carry_f3[1] = 
010101001011110 + 
110101101000000 = 
001010110011110

// TODO: 恢复余数的方法只是自己根据fp64猜的...
msk_dig[2][55:42] = 00000000000010
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[1], 1'b0} | 00000000000010} = 011100111100010
// 111101000000000 + 
// 011100110000000 = 
// 011001110000000

注意, 此时已经求出了12-bit的q
q_real = 1.11001111001
q_real ^ 2 = 11.0100010111010100110001000
a_frac << 1 = 11.0100011000
diff = 0.00000000001010110011110000000

// ======================
rem_sum_in[2] = new_rem_sum_f3[1][14:0] = 010101001011110
rem_carry_in[2] = new_rem_carry_f3[1][14:0] = 110101101000000

rem_sum_msb3[1][5:3] = 010
rem_carry_msb3[1][5:3] = 110
->
quot_dig3[2] = 01
->
prev_quot[2] = new_quot3_f3[1] = 1110011110010
prev_quot_m1[2] = new_quot3_m1_f3[1] = 1110011110000
new_quot3_f3[2] = prev_quot[2] & mask_f3[2][55:43] | msk_dig[2][55:43] = 1110011110011
new_quot3_m1_f3[2] = prev_quot[2] & mask_f3[2][55:43] = 1110011110010


注意, 此时: msk_dig[2][55:43] = 0000000000001, csa_minus_val_sqrt3[2]没有包含msk_dig[2][55:43]的LSB.
所以相当于减数的值变小了
csa_minus_val_sqrt3[2] = {new_quot3_f3[1][11: 1], 1'b0} | msk_dig[2][55:44] = 
110011110010 | 
000000000000 = 
110011110010
csa_minus_val3[2] = {2'b00, csa_minus_val_sqrt3[2]} = 00110011110010
csa_val3[2] = ~csa_minus_val3[2][13:0] = 11001100001101
csa_mux[2][14:0] = {csa_val3[2][13:0], 1'b0} = 110011000011010

rem_sum_in[2][13:0] = 10101001011110
rem_carry_in[2][13:0] = 10101101000000

rem_sum_in[2][13:8] 		= 101010
rem_carry_in[2][13:8] 		= 101011
csa_minus_val3[2][11:8] 	=   1100 -> 0011
rem3_sum_minus[2][5:0] 		= 000010
rem3_carry_minus[2][5:0] 	= 110111
rem_sum_msb3[2][5:0] 		= 000010
rem_carry_msb3[2][5:0] 		= 110111

rem_sum_xor[2][9:0] = 
0010111100 ^ 
1010000000 ^ 
1000011010 = 
0000100110
rem_carry_andor[2][10:0] = 10100110001

new_rem_sum3[2][13:0] = {rem_sum_msb3[2][5:0], rem_sum_xor[2][ 8: 1]} = 00001000010011
new_rem_sum_f3[2] = {new_rem_sum3[2][13: 0], 1'b0} = 000010000100110
new_rem_carry3[2][12:0] = {rem_carry_msb3[2][5:1], rem_carry_andor[2][ 9: 2]} = 1101101001100
new_rem_carry_f3[2] = {new_rem_carry3[2][12: 0], quot_dig3[2][0], 1'b0} = 110110100110010

此时:
new_rem_sum_f3[2] + new_rem_carry_f3[2] = 
000010000100110 + 
110110100110010 = 
111000101011000

010101100111100 - 
010110011110010 = 
111111001001010


按照之前的方法计算的结果:
// TODO: 恢复余数的方法只是自己根据fp64猜的...
下次迭代: msk_dig[0][55:42] = 00000000000001
div_sh[14:0] = {1'b0, {new_quot3_m1_f3[2], 1'b0} | 00000000001000} = 011100111100101
111000101011000 + 
011100111100101 = 
010101100111101

忽略求出的Q的LSB:
div_sh[14:0] = {1'b0, new_quot3_m1_f3[2][12:1], 2'b11} = 011100111100111
111000101011000 + 
011100111100111 = 
010101100111111

rem_sum_plus_d_no_sh[14:0] = new_rem_sum_f3[2][14:0] ^ new_rem_carry_f3[2][14:0] ^ div_sh[14:0] = 
000010000100110 ^ 
110110100110010 ^ 
011100111100111 = 
101000011110011

rem_carry_plus_d_no_sh[14:0] =  {
	  (new_rem_sum_f3[2][13:0] & new_rem_carry_f3[2][13:0])
	| (new_rem_sum_f3[2][13:0] & div_sh[13:0])
	| (new_rem_carry_f3[2][13:0] & div_sh[13:0]),
	1'b0
} = 101101001001100

rem_plus_d_no_sh_xor[14:0] = rem_sum_plus_d_no_sh[14:0] ^ rem_carry_plus_d_no_sh[14:0] = 
101000011110011 ^ 
101101001001100 = 
000101010111111

rem_plus_d_no_sh_or [14:1] = rem_sum_plus_d_no_sh[13:0] | rem_carry_plus_d_no_sh[13:0] = 
01000011110011 | 
01101001001100 = 
01101011111111

000101010111 + 
011010111111 = 
100000010110

101000011110011 + 
101101001001100 = 
010101100111111

问题很多, 还是按照15-bit rem来计算比较方便...


q_real = 1.110011110010
q_real ^ 2 = 11.01000101110101001100010
a_frac << 1 = 11.0100011000
diff = 0.0000000000101011001111000


// ================================================================================================================================================
// iter[4]:
// ================================================================================================================================================
rem_sum_f3[14:0] = 001010111110110
rem_carry_f3[14:0] = 100010000000010

quot_f3[12:0] = 1110011111000
quot_m1_f3[12:0] = 1110011110000

raw_mask_f3 = 11110000000000000
mask_f3[0] = 11111111111110000000000000000000000000000000000000000000
msk_dig[0] = mask_f3[0][55:0] ^ {1'b1, mask_f3[0][55:1]} = 
11111111111110000000000000000000000000000000000000000000 ^ 
11111111111111000000000000000000000000000000000000000000 = 
00000000000001000000000000000000000000000000000000000000
msk_dig_3[0] = msk_dig[0][55:1] | msk_dig[0][54:0] = 
0000000000000100000000000000000000000000000000000000000 |
0000000000001000000000000000000000000000000000000000000 = 
0000000000001100000000000000000000000000000000000000000

mask_f3[1] 		= 11111111111111000000000000000000000000000000000000000000
msk_dig[1] 		= 00000000000000100000000000000000000000000000000000000000
msk_dig_3[1] 	= 0000000000000110000000000000000000000000000000000000000

mask_f3[2] 		= 11111111111111100000000000000000000000000000000000000000
msk_dig[2] 		= 00000000000000010000000000000000000000000000000000000000
msk_dig_3[2] 	= 0000000000000011000000000000000000000000000000000000000



// ================================================================================================================================================
选择常数
0:
m[-1].0 = -13 = 1110_011
m[-0].0 =  -4 = 1111_100
m[+1].0 =  +4 = 0000_100
m[+2].0 = +12 = 0001_100

1:
m[-1].1 = -14 = 1110_010
m[-0].1 =  -5 = 1111_011
m[+1].1 =  +4 = 0000_100
m[+2].1 = +14 = 0001_110

2:
m[-1].2 = -16 = 1110_000
m[-0].2 =  -6 = 1111_010
m[+1].2 =  +4 = 0000_100
m[+2].2 = +16 = 0010_000

3:
m[-1].3 = -17 = 1101_111
m[-0].3 =  -6 = 1111_010
m[+1].3 =  +4 = 0000_100
m[+2].3 = +16 = 0010_000

4:
m[-1].4 = -18 = 1101_110
m[-0].4 =  -6 = 1111_010
m[+1].4 =  +6 = 0000_110
m[+2].4 = +18 = 0010_010

5:
m[-1].5 = -20 = 1101_100
m[-0].5 =  -8 = 1111_000
m[+1].5 =  +6 = 0000_110
m[+2].5 = +20 = 0010_100

6:
m[-1].6 = -22 = 1101_010
m[-0].6 =  -8 = 1111_000
m[+1].6 =  +8 = 0001_000
m[+2].6 = +20 = 0010_100

7:
m[-1].7 = -23 = 1101_001
m[-0].7 =  -8 = 1111_000
m[+1].7 =  +8 = 0001_000
m[+2].7 = +20 = 0010_100

// ================================================================================================================================================
指数是奇数:
a_frac = 1.1010001100
a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
a_frac >> 1 = 0.11010001100
rem[0] = 1 - (a_frac >> 1) = 11_11010001100
s[0] = 1
rt_pos = 01_
rt_neg = 00_
rt[0] = 01_
rt_m[0] = 00_

4 * rem[0] = 1111_01000110000
(4 * rem[0])_trunc_4_3 = 1111_010, belongs to "[m[-0].7, m[+1].7)" -> s[1] = 0
rt_pos  = 01_00
rt_neg  = 00_00
rt[1]   = 01_00
rt_m[1] = 00_11

f[1] = 0
4 * rem[0] + f[1] = 
1111_01000110000 + 
0000_00000000000 = 
1111_01000110000 -> 
rem[1] = 11_01000110000

(4 * rem[1])_trunc_4_3 = 1101_000, belongs to "[-inf, m[-1].7)" -> s[2] = -2
rt_pos  = 01_0000
rt_neg  = 00_0010
rt[2]   = 00_1110
rt_m[2] = 00_1101

f[2] = {rt_m[1] * 4, 11} = 0011_11
4 * rem[1] + f[2] = 
1101_00011000000 + 
0011_11000000000 = 
0000_11011000000 -> 
rem[2] = 00_11011000000

(4 * rem[2])_trunc_4_3 = 0011_011, belongs to "[m[+2].6, +inf)" -> s[3] = +2
rt_pos  = 01_000010
rt_neg  = 00_001000
rt[3]   = 00_111010
rt_m[3] = 00_111001

f[3] = -{(rt[2] * 4).丢弃lsb, 100} = -11_100100
4 * rem[2] + f[3] = 
0011_01100000000 -
0011_10010000000 = 
1111_11010000000 -> 
rem[3] = 11_11010000000


(4 * rem[3])_trunc_4_3 = 1111_010, belongs to "[m[-0].6, m[+1].6)" -> s[4] = 0
rt_pos  = 01_00001000
rt_neg  = 00_00100000
rt[4]   = 00_11101000
rt_m[4] = 00_11100111

f[4] = 0
4 * rem[3] + f[4] = 
1111_010000000000000000000000000000000000 + 
0000_000000000000000000000000000000000000 = 
1111_010000000000000000000000000000000000 -> 
rem[4] = 11_010000000000000000000000000000000000

{(rt_m[4] << 1).丢弃LSB, 1} = 0001_110011101
1111_010000000000000000000000000000000000 + 
0001_110011101000000000000000000000000000 = 
0001_000011101000000000000000000000000000

(4 * rem[4])_trunc_4_3 = 1101_000, belongs to "[-inf, m[-1].6)" -> s[5] = -2
rt_pos  = 01_0000100000
rt_neg  = 00_0010000010
rt[5]   = 00_1110011110
rt_m[5] = 00_1110011101

f[5] = {(rt_m[4] * 4).丢弃低2位, 11} = 0011_10011111
4 * rem[4] + f[5] = 
1101_000000000000000000000000000000000000 + 
0011_100111110000000000000000000000000000 = 
0000_100111110000000000000000000000000000 -> 
rem[5] = 00_100111110000000000000000000000000000

// rem[5] is correct

(4 * rem[5])_trunc_4_3 = 0010_011, belongs to "[m[+1].6, m[+1].6)" -> s[6] = +1
rt_pos  = 01_000010000001
rt_neg  = 00_001000001000
rt[6]   = 00_111001111001
rt_m[6] = 00_111001111000

f[6] = -{rt[5] * 2, 01} = -0001_110011110001
4 * rem[5] + f[6] = 
0010_011111000000000000000000000000000000 -
0001_110011110001000000000000000000000000 = 
0000_101011001111000000000000000000000000 -> 
rem[6] = 00_101011001111000000000000000000000000

// rem[6] is correct

(4 * rem[6])_trunc_4_3 = 0010_101, belongs to "[m[+2].6, +inf)" -> s[7] = +2
rt_pos  = 01_00001000000110
rt_neg  = 00_00100000100000
rt[7]   = 00_11100111100110
rt_m[7] = 00_11100111100101

f[7] = -{(rt[6] * 4).丢弃lsb, 100} = -0011_10011110010100
4 * rem[6] + f[7] = 
0010_101100111100000000000000000000000000 -
0011_100111100101000000000000000000000000 = 
1111_000101010111000000000000000000000000 -> 
rem[7] = 11_000101010111000000000000000000000000

{(rt_m[7] << 1).丢弃LSB, 1} = 01_11001111001011
11_000101010111000000000000000000000000 + 
01_110011110010110000000000000000000000 = 
00_111001001001110000000000000000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.1100111100101
rt_real ^ 2 = 11.010001011111000110110110010
rem_real = 11.0100011000 - 11.010001011111000110110110010 = 
0.00000000000011100100100111000000000000000000000000
// rem[7] is correct

(4 * rem[7])_trunc_4_3 = 1100_010, belongs to "[-inf, m[-1].6)" -> s[8] = -2
rt_pos  = 01_0000100000011000
rt_neg  = 00_0010000010000010
rt[8]   = 00_1110011110010110
rt_m[8] = 00_1110011110010101

f[8] = {(rt_m[7] * 4).丢弃低2位, 11} = 0011_10011110010111
4 * rem[7] + f[8] = 
1100_010101011100000000000000000000000000 +
0011_100111100101110000000000000000000000 = 
1111_111101000001110000000000000000000000 -> 
rem[8] = 11_111101000001110000000000000000000000

{(rt_m[8] << 1).丢弃LSB, 1} = 01_1100111100101011
11_111101000001110000000000000000000000 + 
01_110011110010101100000000000000000000 = 
01_110000110100011100000000000000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.110011110010101
rt_real ^ 2 = 11.010001011111100011110010111001
rem_real = 11.0100011000 - 11.010001011111100011110010111001 = 
0.00000000000001110000110100011100000000000000000000
// rem[8] is correct

(4 * rem[8])_trunc_4_3 = 1111_110, belongs to "[m[-0].6, m[+1].6)" -> s[9] = 0
rt_pos  = 01_000010000001100000
rt_neg  = 00_001000001000001000
rt[9]   = 00_111001111001011000
rt_m[9] = 00_111001111001010111

f[9] = 0
4 * rem[8] + f[9] = 
1111_110100000111000000000000000000000000 +
0000_000000000000000000000000000000000000 = 
1111_110100000111000000000000000000000000 -> 
rem[9] = 11_110100000111000000000000000000000000

{(rt_m[9] << 1).丢弃LSB, 1} = 01_110011110010101111
11_110100000111000000000000000000000000 + 
01_110011110010101111000000000000000000 = 
01_100111111001101111000000000000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.11001111001010111
rt_real ^ 2 = 11.01000101111111100110000001100100010000000000000000
rem_real = 11.0100011000 - 11.01000101111111100110000001100100010000000000000000 = 
0.00000000000000011001111110011011110000000000000000
// rem[9] is correct

(4 * rem[9])_trunc_4_3 = 1111_010, belongs to "[m[-0].6, m[+1].6)" -> s[10] = 0
rt_pos   = 01_00001000000110000000
rt_neg   = 00_00100000100000100000
rt[10]   = 00_11100111100101100000
rt_m[10] = 00_11100111100101011111

f[10] = 0
4 * rem[9] + f[10] = 
1111_010000011100000000000000000000000000 +
0000_000000000000000000000000000000000000 = 
1111_010000011100000000000000000000000000 -> 
rem[10] = 11_010000011100000000000000000000000000

{(rt_m[10] << 1).丢弃LSB, 1} = 01_11001111001010111111
11_010000011100000000000000000000000000 + 
01_110011110010101111110000000000000000 = 
01_000100001110101111110000000000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.1100111100101011111
rt_real ^ 2 = 11.01000101111111111011101111000101000001
rem_real = 11.0100011000 - 11.01000101111111111011101111000101000001 = 
0.00000000000000000100010000111010111111000000000000
// rem[10] is correct

(4 * rem[10])_trunc_4_3 = 1101_000, belongs to "[-inf, m[-1].6)" -> s[11] = -2
rt_pos   = 01_0000100000011000000000
rt_neg   = 00_0010000010000010000010
rt[11]   = 00_1110011110010101111110
rt_m[11] = 00_1110011110010101111101

f[11] = {(rt_m[10] * 4).丢弃低2位, 11} = 0011_10011110010101111111
4 * rem[10] + f[11] = 
1101_000001110000000000000000000000000000 +
0011_100111100101011111110000000000000000 = 
0000_101001010101011111110000000000000000 -> 
rem[11] = 00_101001010101011111110000000000000000


a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.110011110010101111110
rt_real ^ 2 = 11.01000101111111111111010110101010100000010000000000
rem_real = 11.0100011000 - 11.01000101111111111111010110101010100000010000000000 = 
0.00000000000000000000101001010101011111110000000000
// rem[11] is correct

(4 * rem[11])_trunc_4_3 = 0010_100, belongs to "[m[+2].6, +inf)" -> s[12] = +2
rt_pos   = 01_000010000001100000000010
rt_neg   = 00_001000001000001000001000
rt[12]   = 00_111001111001010111111010
rt_m[12] = 00_111001111001010111111001

f[12] = -{(rt[11] * 4).丢弃lsb, 100}= -0011_100111100101011111100100
4 * rem[11] + f[12] = 
0010_100101010101111111000000000000000000 -
0011_100111100101011111100100000000000000 = 
1110_111101110000011111011100000000000000 -> 
rem[12] = 10_111101110000011111011100000000000000

{(rt_m[12] << 1).丢弃LSB, 1} = 01_110011110010101111110011
10_111101110000011111011100000000000000 + 
01_110011110010101111110011000000000000 = 
00_110001100011001111001111000000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.11001111001010111111001
rt_real ^ 2 = 11.01000101111111111111110011100111001100001100010000
rem_real = 11.0100011000 - 11.01000101111111111111110011100111001100001100010000 = 
0.00000000000000000000001100011000110011110011110000
// rem[12] is correct

(4 * rem[12])_trunc_4_3 = 1011_110, belongs to belongs to "[-inf, m[-1].6)" -> s[13] = -2
rt_pos   = 01_00001000000110000000001000
rt_neg   = 00_00100000100000100000100010
rt[13]   = 00_11100111100101011111100110
rt_m[13] = 00_11100111100101011111100101

f[13] = {(rt_m[12] * 4).丢弃低2位, 11} = 0011_100111100101011111100111
4 * rem[12] + f[13] = 
1011_110111000001111101110000000000000000 +
0011_100111100101011111100111000000000000 = 
1111_011110100111011101010111000000000000 -> 
rem[13] = 11_011110100111011101010111000000000000

{(rt_m[13] << 1).丢弃LSB, 1} = 01_11001111001010111111001011
11_011110100111011101010111000000000000 + 
01_110011110010101111110010110000000000 = 
01_010010011010001101001001110000000000

a_frac << 1 = 11.0100011000
sqrt(a_frac << 1) = 1.11001111001010111111001011011011000110001110001001
rt_real = 1.1100111100101011111100101
rt_real ^ 2 = 11.01000101111111111111111010110110010111001011011001
rem_real = 11.0100011000 - 11.01000101111111111111111010110110010111001011011001 = 
0.00000000000000000000000101001001101000110100100111
// rem[13] is correct

此时得到的结果已经足够给f32用来rounding

对于F32来说，迭代6 cycles, 将整数位计算进来，则得到了26-bit结果
如果只要求得到rem[13], 而不需要根据rem[13]得到正确的余数(即在rem[13] < 0时做恢复余数的计算), 那么只需要28-bit的rem和CSA就够了

F64: 迭代13 cycles, 将会得到(13 * 4 + 2) = 54-bit结果, 参考上面, 似乎只需要56-bit就够了, 但是参考论文里用了59-bit
// TODO: 数据通路的宽度还需要测试

// ================================================================================================================================================

指数是奇数:
a_frac = 1.01111111101111111101111
a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
a_frac >> 1 = 0.101111111101111111101111

rem[0] = 1 - (a_frac >> 1) = 11_101111111101111111101111
s[0] = 1
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

(4 * rem[0])_trunc_4_3 = 1110_111, belongs to "[m[-1].7, m[0].7)" -> s[1] = -1
rt_pos  = 01_00
rt_neg  = 00_01
rt[1]   = 00_11
rt_m[1] = 00_10

f[1] = {(rt_m[0] * 2).丢弃最低位, 111} = 0001_11
4 * rem[0] + f[1] = 
1110_111111110111111110111100 + 
0001_110000000000000000000000 = 
0000_101111110111111110111100 -> 
rem[1] = 00_101111110111111110111100

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.1
rt_real ^ 2 = 10.01000000000000000000000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.01000000000000000000000000000000000000000000000000 = 
0.10111111011111111011110000000000000000000000000000
// rem[1] is correct

(4 * rem[1])_trunc_4_3 = 0010_111, belongs to "[m[+2].4, +inf)" -> s[2] = +2
rt_pos  = 01_0010
rt_neg  = 00_0100
rt[2]   = 00_1110
rt_m[2] = 00_1101

f[2] = -{(rt[1] * 4).丢弃lsb, 100}= -0011_0100
4 * rem[1] + f[2] = 
0010_111111011111111011110000 - 
0011_010000000000000000000000 = 
1111_101111011111111011110000 -> 
rem[2] = 11_101111011111111011110000

{(rt_m[2] << 1).丢弃LSB, 1} = 01_1011
11_101111011111111011110000 + 
01_101100000000000000000000 = 
01_011011011111111011110000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.101
rt_real ^ 2 = 10.10100100000000000000000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.10100100000000000000000000000000000000000000000000 = 
0.01011011011111111011110000000000000000000000000000
// rem[2] is correct

(4 * rem[2])_trunc_4_3 = 1110_111, belongs to "[m[-1].6, m[0].6)" -> s[3] = -1
rt_pos  = 01_001000
rt_neg  = 00_010001
rt[3]   = 00_110111
rt_m[3] = 00_110110

f[3] = {(rt_m[2] * 2).丢弃最低位, 111} = 0001_101111
4 * rem[2] + f[3] = 
1110_111101111111101111000000 +
0001_101111000000000000000000 = 
0000_101100111111101111000000 -> 
rem[3] = 00_101100111111101111000000


a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.10111
rt_real ^ 2 = 10.11110100010000000000000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.11110100010000000000000000000000000000000000000000 = 
0.00001011001111111011110000000000000000000000000000
// rem[3] is correct

(4 * rem[3])_trunc_4_3 = 0010_110, belongs to "[m[+2].6, +inf)" -> s[4] = +2
rt_pos  = 01_00100010
rt_neg  = 00_01000100
rt[4]   = 00_11011110
rt_m[4] = 00_11011101

f[4] = -{(rt[3] * 4).丢弃lsb, 100}= -0011_01110100
4 * rem[3] + f[4] = 
0010_110011111110111100000000 -
0011_011101000000000000000000 = 
1111_010110111110111100000000 -> 
rem[4] = 11_010110111110111100000000

{(rt_m[4] << 1).丢弃LSB, 1} = 01_10111011
11_010110111110111100000000 + 
01_101110110000000000000000 = 
01_000101101110111100000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.1011101
rt_real ^ 2 = 10.11111011001001000000000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.11111011001001000000000000000000000000000000000000 = 
0.00000100010110111011110000000000000000000000000000
// rem[4] is correct

(4 * rem[4])_trunc_4_3 = 1101_011, belongs to "[m[-1].6, m[0].6)" -> s[5] = -1
rt_pos  = 01_0010001000
rt_neg  = 00_0100010001
rt[5]   = 00_1101110111
rt_m[5] = 00_1101110110

f[5] = {(rt_m[4] * 2).丢弃最低位, 111} = 0001_1011101111
4 * rem[4] + f[5] = 
1101_011011111011110000000000 +
0001_101110111100000000000000 = 
1111_001010110111110000000000 -> 
rem[5] = 11_001010110111110000000000

{(rt_m[5] << 1).丢弃LSB, 1} = 01_1011101101
11_001010110111110000000000 + 
01_101110110100000000000000 = 
00_111001101011110000000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.101110110
rt_real ^ 2 = 10.11111110100110010000000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.11111110100110010000000000000000000000000000000000 = 
0.00000000111001101011110000000000000000000000000000
// rem[5] is correct

(4 * rem[5])_trunc_4_3 = 1100_101, belongs to "[-inf, m[-1].6)" -> s[6] = -2
rt_pos  = 01_001000100000
rt_neg  = 00_010001000110
rt[6]   = 00_110111011010
rt_m[6] = 00_110111011001

f[6] = {(rt_m[5] * 4).丢弃低2位, 11} = 0011_0111011011
4 * rem[5] + f[6] = 
1100_101011011111000000000000 +
0011_011101101100000000000000 = 
0000_001001001011000000000000 -> 
rem[6] = 00_001001001011000000000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.10111011010
rt_real ^ 2 = 10.11111111011101101001000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011101101001000000000000000000000000000000 = 
0.00000000000010010010110000000000000000000000000000
// rem[6] is correct

(4 * rem[6])_trunc_4_3 = 0000_100, belongs to "[m[-0].6, m[+1].6)" -> s[7] = 0
rt_pos  = 01_00100010000000
rt_neg  = 00_01000100011000
rt[7]   = 00_11011101101000
rt_m[7] = 00_11011101100111

f[7] = 0
4 * rem[6] + f[7] = 
0000_100100101100000000000000 +
0000_000000000000000000000000 = 
0000_100100101100000000000000 -> 
rem[7] = 00_100100101100000000000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.1011101101000
rt_real ^ 2 = 10.11111111011101101001000000000000000000000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011101101001000000000000000000000000000000 = 
0.00000000000010010010110000000000000000000000000000
// rem[7] is correct

(4 * rem[7])_trunc_4_3 = 0010_010, belongs to "[m[+1].6, m[+1].6)" -> s[8] = +1
rt_pos  = 01_0010001000000001
rt_neg  = 00_0100010001100000
rt[8]   = 00_1101110110100001
rt_m[8] = 00_1101110110100000

f[8] = -{rt[7] * 2, 01} = -0001_1011101101000001
4 * rem[7] + f[8] = 
0010_010010110000000000000000 -
0001_101110110100000100000000 = 
0000_100011111011111100000000 -> 
rem[8] = 00_100011111011111100000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.101110110100001
rt_real ^ 2 = 10.11111111011111010111110100000100000000000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011111010111110100000100000000000000000000 = 
0.00000000000000100011111011111100000000000000000000
// rem[8] is correct

(4 * rem[8])_trunc_4_3 = 0010_001, belongs to "[m[+1].6, m[+1].6)" -> s[9] = +1
rt_pos  = 01_001000100000000101
rt_neg  = 00_010001000110000000
rt[9]   = 00_110111011010000101
rt_m[9] = 00_110111011010000100

f[9] = -{rt[8] * 2, 01} = -0001_101110110100001001
4 * rem[8] + f[9] = 
0010_001111101111110000000000 -
0001_101110110100001001000000 = 
0000_100000111011100111000000 -> 
rem[9] = 00_100000111011100111000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.10111011010000101
rt_real ^ 2 = 10.11111111011111110011100001000110010000000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011111110011100001000110010000000000000000 = 
0.00000000000000001000001110111001110000000000000000
// rem[9] is correct

(4 * rem[9])_trunc_4_3 = 0010_000, belongs to "[m[+1].6, m[+1].6)" -> s[10] = +1
rt_pos   = 01_00100010000000010101
rt_neg   = 00_01000100011000000000
rt[10]   = 00_11011101101000010101
rt_m[10] = 00_11011101101000010100

f[10] = -{rt[9] * 2, 01} = -0001_10111011010000101001
4 * rem[9] + f[10] = 
0010_000011101110011100000000 -
0001_101110110100001010010000 = 
0000_010100111010010001110000 -> 
rem[10] = 00_010100111010010001110000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.1011101101000010101
rt_real ^ 2 = 10.11111111011111111010011100010110111001000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011111111010011100010110111001000000000000 = 
0.00000000000000000001010011101001000111000000000000
// rem[10] is correct

(4 * rem[10])_trunc_4_3 = 0001_010, belongs to "[m[+1].6, m[+1].6)" -> s[11] = +1
rt_pos   = 01_0010001000000001010101
rt_neg   = 00_0100010001100000000000
rt[11]   = 00_1101110110100001010101
rt_m[11] = 00_1101110110100001010100

f[11] = -{rt[10] * 2, 01} = -0001_1011101101000010101001
4 * rem[10] + f[11] = 
0001_010011101001000111000000 -
0001_101110110100001010100100 = 
1111_100100110100111100011100 -> 
rem[11] = 11_100100110100111100011100

{(rt_m[11] << 1).丢弃LSB, 1} = 01_1011101101000010101001
11_100100110100111100011100 + 
01_101110110100001010100100 = 
01_010011101001000111000000

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.101110110100001010100
rt_real ^ 2 = 10.11111111011111111010011100010110111001000000000000
rem_real = 10.11111111011111111011110 - 10.11111111011111111010011100010110111001000000000000 = 
0.00000000000000000001010011101001000111000000000000
// rem[11] is correct

(4 * rem[11])_trunc_4_3 = 1110_010, belongs to belongs to "[m[-1].7, m[0].7)" -> s[12] = -1
rt_pos   = 01_001000100000000101010100
rt_neg   = 00_010001000110000000000001
rt[12]   = 00_110111011010000101010011
rt_m[12] = 00_110111011010000101010010

f[12] = {(rt_m[11] * 2).丢弃最低位, 111} = 0001_101110110100001010100111
4 * rem[11] + f[12] = 
1110_010011010011110001110000 +
0001_101110110100001010100111 = 
0000_000010000111111100010111 -> 
rem[12] = 00_000010000111111100010111

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.10111011010000101010011
rt_real ^ 2 = 10.11111111011111111011101111011110000000111010010000
rem_real = 10.11111111011111111011110 - 10.11111111011111111011101111011110000000111010010000 = 
0.00000000000000000000000000100001111111000101110000
// rem[12] is correct

(4 * rem[12])_trunc_4_3 = 0000_001, belongs to belongs to "[m[-0].6, m[+1].6)" -> s[13] = 0
rt_pos   = 01_00100010000000010101010000
rt_neg   = 00_01000100011000000000000100
rt[13]   = 00_11011101101000010101001100
rt_m[13] = 00_11011101101000010101001011

f[13] = 0
4 * rem[12] + f[13] = 
0000_001000011111110001011100 +
0000_000000000000000000000000 = 
0000_001000011111110001011100 -> 
rem[13] = 00_001000011111110001011100

a_frac << 1 = 10.11111111011111111011110
sqrt(a_frac << 1) = 1.10111011010000101010011000001001110100000110010111
rt_real = 1.1011101101000010101001100
rt_real ^ 2 = 10.11111111011111111011101111011110000000111010010000
rem_real = 10.11111111011111111011110 - 10.11111111011111111011101111011110000000111010010000 = 
0.00000000000000000000000000100001111111000101110000
// rem[13] is correct


// ================================================================================================================================================

指数是偶数:
a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
a_frac >> 2 = 0.0111111111100000010111100

rem[0] = 1 - (a_frac >> 2) = 11_0111111111100000010111100
s[0] = 1
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

(4 * rem[0])_trunc_4_3 = 1101_111, belongs to "[m[-1].7, m[0].7)" -> s[1] = -1
rt_pos  = 01_00
rt_neg  = 00_01
rt[1]   = 00_11
rt_m[1] = 00_10

f[1] = {(rt_m[0] * 2).丢弃最低位, 111} = 0001_11
4 * rem[0] + f[1] = 
1101_1111111110000001011110000 + 
0001_1100000000000000000000000 = 
1111_1011111110000001011110000 -> 
rem[1] = 11_1011111110000001011110000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_01
11_1011111110000001011110000 + 
01_0100000000000000000000000 = 
00_1111111110000001011110000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.0
rt_real ^ 2 = 1.00000000000000000000000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.00000000000000000000000000000000000000000000000000 = 
0.11111111100000010111100000000000000000000000000000
// rem[1] is correct

(4 * rem[1])_trunc_4_3 = 1110_111, belongs to "[m[-1].4, m[0].4)" -> s[2] = -1
rt_pos  = 01_0000
rt_neg  = 00_0101
rt[2]   = 00_1011
rt_m[2] = 00_1010

f[2] = {(rt_m[1] * 2).丢弃最低位, 111} = 0001_0111
4 * rem[1] + f[2] = 
1110_1111111000000101111000000 + 
0001_0111000000000000000000000 = 
0000_0110111000000101111000000 -> 
rem[2] = 00_0110111000000101111000000


a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.011
rt_real ^ 2 = 1.11100100000000000000000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11100100000000000000000000000000000000000000000000 = 
0.00011011100000010111100000000000000000000000000000
// rem[2] is correct

(4 * rem[2])_trunc_4_3 = 0001_101, belongs to "[m[+1].3, m[+2].3)" -> s[3] = +1
rt_pos  = 01_000001
rt_neg  = 00_010100
rt[3]   = 00_101101
rt_m[3] = 00_101100

f[3] = -{rt[2] * 2, 01} = -0001_011001
4 * rem[2] + f[3] = 
0001_1011100000010111100000000 -
0001_0110010000000000000000000 = 
0000_0101010000010111100000000 -> 
rem[3] = 00_0101010000010111100000000


a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.01101
rt_real ^ 2 = 1.11111010010000000000000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111010010000000000000000000000000000000000000000 = 
0.00000101010000010111100000000000000000000000000000
// rem[3] is correct

(4 * rem[3])_trunc_4_3 = 0001_010, belongs to "[m[+1].3, m[+2].3)" -> s[4] = +1
rt_pos  = 01_00000101
rt_neg  = 00_01010000
rt[4]   = 00_10110101
rt_m[4] = 00_10110100

f[4] = -{rt[3] * 2, 01} = -0001_01101001
4 * rem[3] + f[4] = 
0001_0101000001011110000000000 -
0001_0110100100000000000000000 = 
1111_1110011101011110000000000 -> 
rem[4] = 11_1110011101011110000000000

{(rt_m[4] << 1).丢弃LSB, 1} = 01_01101001
11_1110011101011110000000000 + 
01_0110100100000000000000000 = 
01_0101000001011110000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.0110100
rt_real ^ 2 = 1.11111010010000000000000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111010010000000000000000000000000000000000000000 = 
0.00000101010000010111100000000000000000000000000000
// rem[4] is correct

(4 * rem[4])_trunc_4_3 = 1111_100, belongs to "[m[0].3, m[+1].3)" -> s[5] = 0
rt_pos  = 01_0000010100
rt_neg  = 00_0101000000
rt[5]   = 00_1011010100
rt_m[5] = 00_1011010011

f[5] = 0
4 * rem[4] + f[5] = 
1111_1001110101111000000000000 +
0000_0000000000000000000000000 = 
1111_1001110101111000000000000 -> 
rem[5] = 11_1001110101111000000000000

{(rt_m[5] << 1).丢弃LSB, 1} = 01_0110100111
11_1001110101111000000000000 + 
01_0110100111000000000000000 = 
01_0000011100111000000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.011010011
rt_real ^ 2 = 1.11111110011110100100000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111110011110100100000000000000000000000000000000 = 
0.00000001000001110011100000000000000000000000000000
// rem[5] is correct

(4 * rem[5])_trunc_4_3 = 1110_011, belongs to "[m[-1].3, m[0].3)" -> s[6] = -1
rt_pos  = 01_000001010000
rt_neg  = 00_010100000001
rt[6]   = 00_101101001111
rt_m[6] = 00_101101001110

f[6] = {(rt_m[5] * 2).丢弃最低位, 111} = 0001_011010011111
4 * rem[5] + f[6] = 
1110_0111010111100000000000000 +
0001_0110100111110000000000000 = 
1111_1101111111010000000000000 -> 
rem[6] = 11_1101111111010000000000000

{(rt_m[6] << 1).丢弃LSB, 1} = 01_011010011101
11_1101111111010000000000000 + 
01_0110100111010000000000000 = 
01_0100100110100000000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.01101001110
rt_real ^ 2 = 1.11111111001011110001000000000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111110011110100100000000000000000000000000000000 = 
0.00000000010100100110100000000000000000000000000000
// rem[6] is correct

(4 * rem[6])_trunc_4_3 = 1111_011, belongs to "[m[0].3, m[+1].3)" -> s[7] = 0
rt_pos  = 01_00000101000000
rt_neg  = 00_01010000000100
rt[7]   = 00_10110100111100
rt_m[7] = 00_10110100111011

f[7] = 0
4 * rem[6] + f[7] = 
1111_0111111101000000000000000 +
0000_0000000000000000000000000 = 
1111_0111111101000000000000000 -> 
rem[7] = 11_0111111101000000000000000

{(rt_m[7] << 1).丢弃LSB, 1} = 01_01101001110111
11_0111111101000000000000000 + 
01_0110100111011100000000000 = 
00_1110100100011100000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.0110100111011
rt_real ^ 2 = 1.11111111011100101110011001000000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111110011110100100000000000000000000000000000000 = 
0.00000000000011101001000111000000000000000000000000
// rem[7] is correct

(4 * rem[7])_trunc_4_3 = 1101_111, belongs to "[m[-1].3, m[0].3)" -> s[8] = -1
rt_pos  = 01_0000010100000000
rt_neg  = 00_0101000000010001
rt[8]   = 00_1011010011101111
rt_m[8] = 00_1011010011101110

f[8] = {(rt_m[7] * 2).丢弃最低位, 111} = 0001_0110100111011111
4 * rem[7] + f[8] = 
1101_1111110100000000000000000 +
0001_0110100111011111000000000 = 
1111_0110011011011111000000000 -> 
rem[8] = 11_0110011011011111000000000

{(rt_m[8] << 1).丢弃LSB, 1} = 01_0110100111011101
11_0110011011011111000000000 + 
01_0110100111011101000000000 = 
00_1101000010111100000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.011010011101110
rt_real ^ 2 = 1.11111111011111100011010100010000000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111111011111100011010100010000000000000000000000 = 
0.00000000000000110100001011110000000000000000000000
// rem[8] is correct

(4 * rem[8])_trunc_4_3 = 1101_100, belongs to "[-inf, m[-1].3)" -> s[9] = -2
rt_pos  = 01_000001010000000000
rt_neg  = 00_010100000001000110
rt[9]   = 00_101101001110111010
rt_m[9] = 00_101101001110111001

f[9] = {(rt_m[8] * 4).丢弃低2位, 11} = 0010_1101001110111011
4 * rem[8] + f[9] = 
1101_1001101101111100000000000 +
0010_1101001110111011000000000 = 
0000_0110111100110111000000000 -> 
rem[9] = 00_0110111100110111000000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.01101001110111010
rt_real ^ 2 = 1.11111111100000010000100011001001000000000000000000
rem_real = 1.11111111100000010111100 - 1.11111111100000010000100011001001000000000000000000 = 
0.00000000000000000110111100110111000000000000000000
// rem[9] is correct

(4 * rem[9])_trunc_4_3 = 0001_101, belongs to "[m[+1].3, m[+2].3)" -> s[10] = +1
rt_pos   = 01_00000101000000000001
rt_neg   = 00_01010000000100011000
rt[10]   = 00_10110100111011101001
rt_m[10] = 00_10110100111011101000

f[10] = -{rt[9] * 2, 01} = -0001_01101001110111010001
4 * rem[9] + f[10] = 
0001_1011110011011100000000000 -
0001_0110100111011101000100000 = 
0000_0101001011111110111100000 -> 
rem[10] = 00_0101001011111110111100000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.0110100111011101001
rt_real ^ 2 = 1.11111111100000010110001101000000010001000000000000
rem_real = 1.11111111100000010111100 - 1.11111111100000010110001101000000010001000000000000 = 
0.00000000000000000001010010111111101111000000000000
// rem[10] is correct

(4 * rem[10])_trunc_4_3 = 0001_010, belongs to "[m[+1].3, m[+2].3)" -> s[11] = +1
rt_pos   = 01_0000010100000000000101
rt_neg   = 00_0101000000010001100000
rt[11]   = 00_1011010011101110100101
rt_m[11] = 00_1011010011101110100100

f[11] = -{rt[10] * 2, 01} = -0001_0110100111011101001001
4 * rem[10] + f[11] = 
0001_0100101111111011110000000 -
0001_0110100111011101001001000 = 
1111_1110001000011110100111000 -> 
rem[11] = 11_1110001000011110100111000

{(rt_m[11] << 1).丢弃LSB, 1} = 01_0110100111011101001001
11_1110001000011110100111000 + 
01_0110100111011101001001000 = 
01_0100101111111011110000000

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.011010011101110100100
rt_real ^ 2 = 1.11111111100000010110001101000000010001000000000000
rem_real = 1.11111111100000010111100 - 1.11111111100000010110001101000000010001000000000000 = 
0.00000000000000000001010010111111101111000000000000
// rem[11] is correct

(4 * rem[11])_trunc_4_3 = 1111_100, belongs to "[m[0].3, m[+1].3)" -> s[12] = 0
rt_pos   = 01_000001010000000000010100
rt_neg   = 00_010100000001000110000000
rt[12]   = 00_101101001110111010010100
rt_m[12] = 00_101101001110111010010011

f[12] = 0
4 * rem[11] + f[12] = 
1111_1000100001111010011100000 +
0000_0000000000000000000000000 = 
1111_1000100001111010011100000 -> 
rem[12] = 11_1000100001111010011100000

{(rt_m[12] << 1).丢弃LSB, 1} = 01_011010011101110100100111
11_1000100001111010011100000 + 
01_0110100111011101001001110 = 
00_1111001001010111100101110

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.01101001110111010010011
rt_real ^ 2 = 1.11111111100000010111010000110110101000011010010000
rem_real = 1.11111111100000010111100 - 1.11111111100000010111010000110110101000011010010000 = 
0.00000000000000000000001111001001010111100101110000
// rem[12] is correct

(4 * rem[12])_trunc_4_3 = 1110_001, belongs to "[m[-1].3, m[0].3)" -> s[13] = -1
rt_pos   = 01_00000101000000000001010000
rt_neg   = 00_01010000000100011000000001
rt[13]   = 00_10110100111011101001001111
rt_m[13] = 00_10110100111011101001001110

0001_01101001110111010010011111
f[13] = {(rt_m[12] * 2).丢弃最低位, 111} = 0001_01101001110111010010011111
4 * rem[12] + f[13] = 
1110_00100001111010011100000000 +
0001_01101001110111010010011111 = 
1111_10001011110001101110011111 -> 
rem[13] = 11_10001011110001101110011111

其实这里就可以停止了...

{(rt_m[13] << 1).丢弃LSB, 1} = 01_01101001110111010010011101
11_10001011110001101110011111 + 
01_01101001110111010010011101 = 
00_11110101101001000000111100

a_frac = 1.11111111100000010111100
sqrt(a_frac) = 1.01101001110111010010011101010110111000111001110010
rt_real = 1.0110100111011101001001110
rt_real ^ 2 = 1.11111111100000010111011100001010010110111111000100
rem_real = 1.11111111100000010111100 - 1.11111111100000010111011100001010010110111111000100 = 
0.00000000000000000000000011110101101001000000111100
// rem[13] is correct


// ================================================================================================================================================
F16: 迭代3个cycles, 迭代完成时得到14位小数，按照上面的分析，应该需要16-bit的rem和csa
指数是偶数:
a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
a_frac >> 2 = 0.011100111101

尝试用rem_s, rem_c的高8位来QDS

rem[0] = 1 - (a_frac >> 2) = 11_01110011110100
rem_s[0] = 1101110011110100
rem_c[0] = 0000000000000000
s[0] = 1
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

(4 * rem[0])_trunc_4_3 = 1101_110, belongs to "[m[-1].7, m[0].7)" -> s[1] = -1
rt_pos  = 01_00
rt_neg  = 00_01
rt[1]   = 00_11
rt_m[1] = 00_10
(rem_s[0][MSB -: 8] + rem_c[0][MSB -: 8]) * 4 = 
11011100 + 
00000000 = 
1101_1100, belongs to "[m[-1].7, m[0].7)" -> s[1] = -1


f[1] = {(rt_m[0] * 2).丢弃最低位, 111} = 0001_11
4 * rem[0] + f[1] = 
1101_11001111010000 + 
0001_11000000000000 = 
1111_10001111010000 -> 
rem[1] = 11_10001111010000
ren_s[1] = 0111001111010000
ren_c[1] = 0111000000000000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_01
11_10001111010000 + 
01_01000000000000 = 
00_11001111010000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.0
rt_real ^ 2 = 1.00000000000000000000000000000000000000000000000000
rem_real = 1.1100111101 - 1.00000000000000000000000000000000000000000000000000 = 
0.11001111010000000000000000000000000000000000000000
// rem[1] is correct

(4 * rem[1])_trunc_4_3 = 1110_001, belongs to "[m[-1].3, m[0].3)" -> s[2] = -1
rt_pos  = 01_0000
rt_neg  = 00_0101
rt[2]   = 00_1011
rt_m[2] = 00_1010
(rem_s[0][MSB -: 8] + rem_c[0][MSB -: 8]) * 4 = 
01110011 + 
01110000 = 
1110_0011, belongs to "[m[-1].3, m[0].3)" -> s[2] = -1

f[2] = {(rt_m[1] * 2).丢弃最低位, 111} = 0001_0111
4 * rem[1] + f[2] = 
1110_00111101000000 + 
0001_01110000000000 = 
1111_10101101000000 -> 
rem[2] = 11_10101101000000
ren_s[2] = 0101001101000000
ren_c[2] = 1001100000000000

{(rt_m[2] << 1).丢弃LSB, 1} = 01_0101
11_10101101000000 + 
01_01010000000000 = 
00_11111101000000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.010
rt_real ^ 2 = 1.10010000000000000000000000000000000000000000000000
rem_real = 1.1100111101 - 1.10010000000000000000000000000000000000000000000000 = 
0.00111111010000000000000000000000000000000000000000
// rem[2] is correct

(4 * rem[2])_trunc_4_3 = 1110_101, belongs to "[m[-1].2, m[0].2)" -> s[3] = -1
rt_pos  = 01_000000
rt_neg  = 00_010101
rt[3]   = 00_101011
rt_m[3] = 00_101010
(rem_s[2][MSB -: 8] + rem_c[2][MSB -: 8]) * 4 = 
01010011 + 
10011000 = 
1110_1011, belongs to "[m[-1].2, m[0].2)" -> s[3] = -1

f[3] = {(rt_m[2] * 2).丢弃最低位, 111} = 0001_010111
4 * rem[2] + f[3] = 
1110_10110100000000 + 
0001_01011100000000 = 
0000_00010000000000 -> 
rem[3] = 00_00010000000000
ren_s[3] = 0111101000000000
ren_c[3] = 1000101000000000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.01011
rt_real ^ 2 = 1.11001110010000000000000000000000000000000000000000
rem_real = 1.1100111101 - 1.11001110010000000000000000000000000000000000000000 = 
0.00000001000000000000000000000000000000000000000000
// rem[3] is correct

(4 * rem[3])_trunc_4_3 = 0000_010, belongs to "[m[0].2, m[+1].2)" -> s[4] = 0
rt_pos  = 01_00000000
rt_neg  = 00_01010100
rt[4]   = 00_10101100
rt_m[4] = 00_10101011
(rem_s[3][MSB -: 8] + rem_c[3][MSB -: 8]) * 4 = 
01111010 + 
10001010 = 
0000_0100, belongs to "[m[0].2, m[+1].2)" -> s[4] = 0

f[4] = 0
4 * rem[3] + f[4] = 
0000_01000000000000 + 
0000_00000000000000 = 
0000_01000000000000 -> 
rem[4] = 00_01000000000000
ren_s[4] = 1110100000000000
ren_c[4] = 0010100000000000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.0101100
rt_real ^ 2 = 1.11001110010000000000000000000000000000000000000000
rem_real = 1.1100111101 - 1.11001110010000000000000000000000000000000000000000 = 
0.00000001000000000000000000000000000000000000000000
// rem[4] is correct

(4 * rem[4])_trunc_4_3 = 0001_000, belongs to "[m[+1].2, m[+2].2)" -> s[5] = +1
rt_pos  = 01_0000000001
rt_neg  = 00_0101010000
rt[5]   = 00_1010110001
rt_m[5] = 00_1010110000
(rem_s[4][MSB -: 8] + rem_c[4][MSB -: 8]) * 4 = 
11101000 + 
00101000 = 
0001_0000, belongs to "[m[+1].2, m[+2].2)" -> s[5] = +1

f[5] = -{rt[4] * 2, 01} = -0001_0101100001
4 * rem[4] + f[5] = 
0001_00000000000000 -
0001_01011000010000 = 
1111_10100111110000 -> 
rem[5] = 11_10100111110000
ren_s[5] = 1010100111101111
ren_c[5] = 0100000000000001

{(rt_m[5] << 1).丢弃LSB, 1} = 01_0101100001
11_10100111110000 + 
01_01011000010000 = 
01_00000000000000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.010110000
rt_real ^ 2 = 1.11001110010000000000000000000000000000000000000000
rem_real = 1.1100111101 - 1.11001110010000000000000000000000000000000000000000 = 
0.00000001000000000000000000000000000000000000000000
// rem[5] is correct

(4 * rem[5])_trunc_4_3 = 1110_100, belongs to "[m[-1].2, m[0].2)" -> s[6] = -1
rt_pos  = 01_000000000100
rt_neg  = 00_010101000001
rt[6]   = 00_101011000011
rt_m[6] = 00_101011000010
(rem_s[5][MSB -: 8] + rem_c[5][MSB -: 8]) * 4 = 
10101001 + 
01000000 = 
1110_1001, belongs to "[m[-1].2, m[0].2)" -> s[6] = -1

f[6] = {(rt_m[5] * 2).丢弃最低位, 111} = 0001_010110000111
4 * rem[5] + f[6] = 
1110_10011111000000 +
0001_01011000011100 = 
1111_11110111011100 -> 
rem[6] = 11_11110111011100
ren_s[6] = 1111000110100100
ren_c[6] = 0000110000111000

{(rt_m[6] << 1).丢弃LSB, 1} = 01_010110000101
11_11110111011100 + 
01_01011000010100 = 
01_01001111110000

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.01011000010
rt_real ^ 2 = 1.11001110111011000001000000000000000000000000000000
rem_real = 1.1100111101 - 1.11001110111011000001000000000000000000000000000000 = 
0.00000000010100111111000000000000000000000000000000
// rem[6] is correct

(4 * rem[6])_trunc_4_3 = 1111_110, belongs to "[m[0].2, m[+1].2)" -> s[7] = 0
rt_pos  = 01_00000000010000
rt_neg  = 00_01010100000100
rt[7]   = 00_10101100001100
rt_m[7] = 00_10101100001011
(rem_s[6][MSB -: 8] + rem_c[6][MSB -: 8]) * 4 = 
11110001 + 
00001100 = 
1111_1101, belongs to "[m[0].2, m[+1].2)" -> s[7] = 0

f[7] = 0
4 * rem[6] + f[7] = 
1111_11011101110000 +
0000_00000000000000 = 
1111_11011101110000 -> 
rem[7] = 11_11011101110000

{(rt_m[7] << 1).丢弃LSB, 1} = 01_01011000010111
11_11011101110000 + 
01_01011000010111 = 
01_00110110000111

a_frac = 1.1100111101
sqrt(a_frac) = 1.01011000010111110011010001010000011010111100010001
rt_real = 1.0101100001011
rt_real ^ 2 = 1.11001111001011001001111001000000000000000000000000
rem_real = 1.1100111101 - 1.11001111001011001001111001000000000000000000000000 = 
0.00000000000100110110000111000000000000000000000000
// rem[7] is correct


// ================================================================================================================================================
F16: 迭代3个cycles, 迭代完成时得到14位小数，按照上面的分析，应该需要16-bit的rem和csa
指数是奇数:
a_frac = 1.1101100111
a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
a_frac >> 1 = 0.11101100111

rem[0] = 1 - (a_frac >> 1) = 11_11101100111000
s[0] = 1
rt_pos  = 01_
rt_neg  = 00_
rt[0]   = 01_
rt_m[0] = 00_

(4 * rem[0])_trunc_4_3 = 1111_101, belongs to "[m[0].7, m[+1].7)" -> s[1] = 0
rt_pos  = 01_00
rt_neg  = 00_00
rt[1]   = 01_00
rt_m[1] = 00_11

f[1] = 0
4 * rem[0] + f[1] = 
1111_10110011100000 + 
0000_00000000000000 = 
1111_10110011100000 -> 
rem[1] = 11_10110011100000

{(rt_m[1] << 1).丢弃LSB, 1} = 01_11
11_10110011100000 + 
01_11000000000000 = 
01_01110011100000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.1
rt_real ^ 2 = 10.01000000000000000000000000000000000000000000000000
rem_real = 11.1011001110 - 10.01000000000000000000000000000000000000000000000000 = 
1.01110011100000000000000000000000000000000000000000
// rem[1] is correct

(4 * rem[1])_trunc_4_3 = 1110_110, belongs to "[m[-1].7, m[0].7)" -> s[2] = -1
rt_pos  = 01_0000
rt_neg  = 00_0001
rt[2]   = 00_1111
rt_m[2] = 00_1110

f[2] = {(rt_m[1] * 2).丢弃最低位, 111} = 0001_1111
4 * rem[1] + f[2] = 
1110_11001110000000 + 
0001_11110000000000 = 
0000_10111110000000 -> 
rem[2] = 00_10111110000000


a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.111
rt_real ^ 2 = 11.10000100000000000000000000000000000000000000000000
rem_real = 11.1011001110 - 11.10000100000000000000000000000000000000000000000000 = 
0.00101111100000000000000000000000000000000000000000
// rem[2] is correct

(4 * rem[2])_trunc_4_3 = 0010_111, belongs to "[m[+2].7, +inf)" -> s[3] = +2
rt_pos  = 01_000010
rt_neg  = 00_000100
rt[3]   = 00_111110
rt_m[3] = 00_111101

f[3] = -{(rt[2] * 4).丢弃lsb, 100}= -0011_110100
4 * rem[2] + f[3] = 
0010_11111000000000 -
0011_11010000000000 = 
1111_00101000000000 -> 
rem[3] = 11_00101000000000

{(rt_m[3] << 1).丢弃LSB, 1} = 01_111011
11_00101000000000 + 
01_11101100000000 = 
01_00010100000000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.11101
rt_real ^ 2 = 11.10100010010000000000000000000000000000000000000000
rem_real = 11.1011001110 - 11.10100010010000000000000000000000000000000000000000 = 
0.00010001010000000000000000000000000000000000000000
// rem[3] is correct

(4 * rem[3])_trunc_4_3 = 1100_101, belongs to "[-inf, m[-1].7)" -> s[4] = -2
rt_pos  = 01_00001000
rt_neg  = 00_00010010
rt[4]   = 00_11110110
rt_m[4] = 00_11110101

f[4] = {(rt_m[3] * 4).丢弃低2位, 11} = 0011_110111
4 * rem[3] + f[4] = 
1100_10100000000000 +
0011_11011100000000 = 
0000_01111100000000 -> 
rem[4] = 00_01111100000000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.1110110
rt_real ^ 2 = 11.10110001100100000000000000000000000000000000000000
rem_real = 11.1011001110 - 11.10110001100100000000000000000000000000000000000000 = 
0.00000001111100000000000000000000000000000000000000
// rem[4] is correct

(4 * rem[4])_trunc_4_3 = 0001_111, belongs to "[m[+1].7, m[+2].7)" -> s[5] = +1
rt_pos  = 01_0000100001
rt_neg  = 00_0001001000
rt[5]   = 00_1111011001
rt_m[5] = 00_1111011000

f[5] = -{rt[4] * 2, 01} = -0001_1110110001
4 * rem[4] + f[5] = 
0001_11110000000000 -
0001_11101100010000 = 
0000_00000011110000 -> 
rem[5] = 00_00000011110000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.111011001
rt_real ^ 2 = 11.10110011011111000100000000000000000000000000000000
rem_real = 11.1011001110 - 11.10110011011111000100000000000000000000000000000000 = 
0.00000000000000111100000000000000000000000000000000
// rem[5] is correct

(4 * rem[5])_trunc_4_3 = 0000_000, belongs to "[m[0].7, m[+1].7)" -> s[6] = 0
rt_pos  = 01_000010000100
rt_neg  = 00_000100100000
rt[6]   = 00_111101100100
rt_m[6] = 00_111101100011

f[6] = 0
4 * rem[5] + f[6] = 
0000_00001111000000 +
0000_00000000000000 = 
0000_00001111000000 -> 
rem[6] = 00_00001111000000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.11101100100
rt_real ^ 2 = 11.10110011011111000100000000000000000000000000000000
rem_real = 11.1011001110 - 11.10110011011111000100000000000000000000000000000000 = 
0.00000000000000111100000000000000000000000000000000
// rem[6] is correct

(4 * rem[6])_trunc_4_3 = 0000_001, belongs to "[m[0].7, m[+1].7)" -> s[7] = 0
rt_pos  = 01_00001000010000
rt_neg  = 00_00010010000000
rt[7]   = 00_11110110010000
rt_m[7] = 00_11110110001111

f[7] = 0
4 * rem[6] + f[7] = 
0000_00111100000000 +
0000_00000000000000 = 
0000_00111100000000 -> 
rem[7] = 00_00111100000000

a_frac << 1 = 11.1011001110
sqrt(a_frac << 1) = 1.11101100100000001111100110000000011001110010001011
rt_real = 1.1110110010000
rt_real ^ 2 = 11.10110011011111000100000000000000000000000000000000
rem_real = 11.1011001110 - 11.10110011011111000100000000000000000000000000000000 = 
0.00000000000000111100000000000000000000000000000000
// rem[7] is correct







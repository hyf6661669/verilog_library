接"test_0.sv", 测试一下参考文献是否能准确求出余数。
选择函数来自于参考论文的"Fig. 6 (c)":
case(w_sum[i][MSB-1:MSB-2], w_carry[i][MSB-1:MSB-2])
	4'b00_00:	q[i+1] = +1;
	4'b00_01:	q[i+1] = +1;
	4'b00_10:	q[i+1] = +0;
	4'b00_11:	q[i+1] = +0;
	4'b01_00:	q[i+1] = +1;
	4'b01_01:	q[i+1] = +2;
	4'b01_10:	q[i+1] = +0;
	4'b01_11:	q[i+1] = +0;
	4'b10_00:	q[i+1] = -0;
	4'b10_01:	q[i+1] = -0;
	4'b10_10:	q[i+1] = -2;
	4'b10_11:	q[i+1] = -1;
	4'b11_00:	q[i+1] = -0;
	4'b11_01:	q[i+1] = -0;
	4'b11_10:	q[i+1] = -1;
	4'b11_11:	q[i+1] = -1;
endcase

// ---------------------------------------------------------------------------------------------------------------------------------------
根据论文对其算法的属性的描述，以及从下面的例子可以得到如下结论:
设最后一次迭代产生的商为Q[n], 对应的部分余数为W[n] = w[n] / 2, 商的绝对值为"quotient", 规格化之前的余数为"remainder", 则有4种情况:
1. W[n]属于区间"[+ D, +2D)" -> quotient = Q[n] + 1, remainder = W[n] - D;
2. W[n]属于区间"[+ 0, + D)" -> quotient = Q[n], remainder = W[n];
3. W[n]属于区间"[- D, - 0)" -> quotient = Q[n] - 1, remainder = W[n] + D;
4. W[n]属于区间"[-2D, - D)" -> quotient = Q[n] - 2, remainder = W[n] + 2D;
总的来说, 至少需要7个全加计算:
fa[0] = w_sum + w_carry;
fa[1] = fa[0] + (-D);
fa[2] = fa[0] + D;
fa[3] = fa[0] + 2D;
fa[4] = Q[n] + 1;
fa[5] = Q[n] - 1;
fa[6] = Q[n] - 2;

在标准的SRT算法中:
rem = rem_sum + rem_carry
rem属于区间"[-D, +D)".
这就导致这个算法在做后处理的时候会比较困难..
为了知道到底应该如何对quotient和remainder进行调整，理论上需要先使用"full-width"的"CPA"将W[n]算出来之后, 再将其和"-D/+D"的大小进行对比。
实际上"fa[0], fa[1], fa[2]"的计算可以是并行的, 但是这么多"full adder"的开销也挺大的, 想办法和前处理步骤中用来求绝对值的全加器复用。
// ---------------------------------------------------------------------------------------------------------------------------------------


先考察简单点的情况:
WIDTH = 24;

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000000010101011 = 171
Q[WIDTH-1:0] = X / D = 4193 = 000000000001000001100001
REM[WIDTH-1:0] = 717047 - 171 * 4193 = 44 = 000000000000000000101100

CLZ_X = 4
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 12
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 14
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101011110000111101110000
Divisor[WIDTH-1:0] 		= 101010110000000000000000

+ D[(WIDTH + 2)-1:0] = 001_01010110000000000000000
+2D[(WIDTH + 2)-1:0] = 010_10101100000000000000000
- D[(WIDTH + 2)-1:0] = 110_10101010000000000000000
-2D[(WIDTH + 2)-1:0] = 101_01010100000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[14];
w[final] = 001_01100000000000000000000 >= 0
// 最后一次迭代的商
q[14] = 0
q_pos = 1000_0100_0000_00
q_neg = 0000_0000_1111_10
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
0010000011000010
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 001000001100001
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
001011000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
001011000000000000000000 >> 16 = 
000000000000000000101100

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 2)-1:0] =  001_01011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0


// 前处理过程中的优化
w_sum_translation[0][WIDTH-1] = Dividend[WIDTH-1] = 1'b1, ~D[WIDTH-1] = ~Divisor[WIDTH-1] = 1'b0, 因此必然有:
w_sum_translation[1][WIDTH] = 1'b1;
w_sum_translation[1][WIDTH-1] = Dividend[WIDTH-2] ^ ~Divisor[WIDTH-2];
w_carry_translation[1][WIDTH] = Dividend[WIDTH-2] & ~Divisor[WIDTH-2];
w_carry_translation[1][WIDTH-1] = Dividend[WIDTH-3] & ~Divisor[WIDTH-3];
按照商选择函数的定义, w_sum_translation[1][WIDTH] = 1'b1, 则q[2]只能是0/-1/-2, 那么就可以快速的根据3-bit信号:
{w_sum_translation[1][WIDTH-1], w_carry_translation[1][WIDTH:WIDTH-1]}
快速确定"q[2]", 从而可以算出:
w_sum_translation[2]
w_carry_translation[2]
由{w_sum_translation[1][WIDTH-1], w_carry_translation[1][WIDTH:WIDTH-1]}的表达式可知, 进一步的, 可以使用4-bit信号:
{Dividend[WIDTH-2:WIDTH-3], Divisor[WIDTH-2:WIDTH-3]}
快速确定"q[2]".
这样相当于补偿了此算法相比于标准"Radix-2 SRT"算法需要的多一次迭代.

比如在这个例子中:
~D[(WIDTH + 2)-1:0] = 110_10101001111111111111111
w_sum_translation[1] = 2 * (w[0] ^ ~D) = 
001_01011110000111101110000 ^ 110_10101001111111111111111 = 
111_11101111110000100011110
w_carry_translation[1] = 2 * (csa_carry(w_sum_translation[0], 0, ~D) | 1'b1) = 
2 * 000_00010000001111011100001 = 
000_00100000011110111000010

加入上述优化之后，意味着前处理过程中需要求出{w_sum_translation[2], w_carry_translation[2]}, 大概会引入:
1. 3-2 CSA的延时.
2. Paper中描述的"Doubling And Translation"所需的延时.
理论分析来看这个延时还是比较小的, 应该不会对Timing造成什么压力.


// 规格化之后必然有:
// q[1] = 1
// 为了方便人工计算，在草稿中一般可以直接令w_carry[1] = -2D, 实际的RTL实现中，是不知道-2D的值的(因为需要对D进行取反，然后再进行一个WIDTH宽度的全加操作).
w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
111_11101000001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_00101000000000000000000
w_sum_translation[1] = 111_11101000001111011100000
w_carry_translation[1] = 000_00101000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_00 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01011110000111101110000 +
	110_10101010000000000000000
) = 2 * 000_00001000000111101110000 = 
000_00010000001111011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11010000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_01010000000000000000000
w_sum_translation[2] = 111_11010000011110111000000
w_carry_translation[2] = 000_01010000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 11_00 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_00010000001111011100000 +
	000_00000000000000000000000
) = 2 * 000_00010000001111011100000 = 
000_00100000011110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_10100000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_10100000000000000000000
w_sum_translation[3] = 111_10100000111101110000000
w_carry_translation[3] = 000_10100000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_00 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00100000011110111000000 +
	000_00000000000000000000000
) = 2 * 000_00100000011110111000000 = 
000_01000000111101110000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_01000001111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_01000000000000000000000
w_sum_translation[4] = 111_01000001111011100000000
w_carry_translation[4] = 001_01000000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_01 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_01000000111101110000000 +
	000_00000000000000000000000
) = 2 * 000_01000000111101110000000 = 
000_10000001111011100000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_10000011110111000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
010_10000000000000000000000
w_sum_translation[5] = 000_10000011110111000000000
w_carry_translation[5] = 000_10000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_00 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_10000001111011100000000 +
	000_00000000000000000000000
) = 2 * 000_10000001111011100000000 = 
001_00000011110111000000000
q_pos = 1000_01
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_01010011101110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
110_00001000000000000000000
w_sum_translation[6] = 001_01010011101110000000000
w_carry_translation[6] = 110_00001000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	001_00000011110111000000000 +
	110_10101010000000000000000
) = 2 * 111_10101101110111000000000 = 
111_01011011101110000000000
q_pos = 1000_010
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_10100111011100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
100_00010000000000000000000
w_sum_translation[7] = 000_10100111011100000000000
w_carry_translation[7] = 110_00010000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_10 -> q[8] = 0
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	111_01011011101110000000000 +
	000_00000000000000000000000
) = 2 * 111_01011011101110000000000 = 
110_10110111011100000000000
q_pos = 1000_0100
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
001_01001110111000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
100_00100000000000000000000
w_sum_translation[8] = 111_01001110111000000000000
w_carry_translation[8] = 110_00100000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 11_10 -> q[9] = -1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	110_10110111011100000000000 +
	000_00000000000000000000000
) = 2 * 110_10110111011100000000000 = 
101_01101110111000000000000
q_pos = 1000_0100_0
q_neg = 0000_0000_1

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
100_01110001110000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
001_00011000000000000000000
w_sum_translation[9] = 110_01110001110000000000000
w_carry_translation[9] = 111_00011000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_11 -> q[10] = -1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	101_01101110111000000000000 +
	001_01010110000000000000000
) = 2 * 110_11000100111000000000000 = 
101_10001001110000000000000
q_pos = 1000_0100_00
q_neg = 0000_0000_11

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
100_01111111100000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_01000000000000000000000
w_sum_translation[10] = 110_01111111100000000000000
w_carry_translation[10] = 111_01000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 10_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	101_10001001110000000000000 +
	001_01010110000000000000000
) = 2 * 110_11011111110000000000000 = 
101_10111111100000000000000
q_pos = 1000_0100_000
q_neg = 0000_0000_111

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_11010011000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
001_01011000000000000000000
w_sum_translation[11] = 110_11010011000000000000000
w_carry_translation[11] = 111_01011000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_11 -> q[12] = -1
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	101_10111111100000000000000 +
	001_01010110000000000000000
) = 2 * 111_00010101100000000000000 = 
110_00101011000000000000000
q_pos = 1000_0100_0000
q_neg = 0000_0000_1111

w_sum[12] = 2 * csa_sum(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
101_10111010000000000000000
w_carry[12] = 2 * csa_carry(w_sum_translation[11], w_carry_translation[11], -q[12] * D) = 
001_01001000000000000000000
w_sum_translation[12] = 111_10111010000000000000000
w_carry_translation[12] = 111_01001000000000000000000
{w_sum_translation[12][MSB-1:MSB-2], w_carry_translation[12][MSB-1:MSB-2]} = 11_11 -> q[13] = -1
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	110_00101011000000000000000 +
	001_01010110000000000000000
) = 2 * 111_10000001000000000000000 = 
111_00000010000000000000000
q_pos = 1000_0100_0000_0
q_neg = 0000_0000_1111_1

w_sum[13] = 2 * csa_sum(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
111_01001000000000000000000
w_carry[13] = 2 * csa_carry(w_sum_translation[12], w_carry_translation[12], -q[13] * D) = 
001_01101000000000000000000
w_sum_translation[13] = 111_01001000000000000000000
w_carry_translation[13] = 001_01101000000000000000000
{w_sum_translation[13][MSB-1:MSB-2], w_carry_translation[13][MSB-1:MSB-2]} = 11_01 -> q[14] = 0
w[13] = 2 * (w[12] - q[13] * D) = 2 * (
	111_00000010000000000000000 +
	001_01010110000000000000000
) = 2 * 000_01011000000000000000000 = 
000_10110000000000000000000
q_pos = 1000_0100_0000_00
q_neg = 0000_0000_1111_10

// 求出最后一次迭代的余数
w[14] = 2 * (w[13] - q[14] * D) = 2 * (
	000_10110000000000000000000 +
	000_00000000000000000000000
) = 2 * 000_10110000000000000000000 = 
001_01100000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000010110010111011 = 11451
Q[WIDTH-1:0] = X / D = 62 = 000000000000000000111110
REM[WIDTH-1:0] = 717047 - 11451 * 62 = 7085 = 000000000001101110101101

CLZ_X = 4
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 6
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 8
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101011110000111101110000
Divisor[WIDTH-1:0] 		= 101100101110110000000000

+ D[(WIDTH + 2)-1:0] = 001_01100101110110000000000
+2D[(WIDTH + 2)-1:0] = 010_11001011101100000000000
- D[(WIDTH + 2)-1:0] = 110_10011010001010000000000
-2D[(WIDTH + 2)-1:0] = 101_00110100010100000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8];
w[final] = 101_11011110010000000000000 < 0
// 最后一次迭代的商
q[8] = 0
q_pos = 1000_0110
q_neg = 0000_1000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
01111101
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0111110
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1_01110111100100000000000 + 1_01100101110110000000000 = 
011011101011010000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
011011101011010000000000 >> 10 = 
000000000001101110101101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_01011110000111101110000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

// 规格化之后必然有:
// q[1] = 1
// 为了方便人工计算，在草稿中一般可以直接令w_carry[1] = -2D, 实际的RTL实现中，是不知道-2D的值的(因为需要对D进行取反，然后再进行一个WIDTH宽度的全加操作).
w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_10111100001111011100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_00110100010100000000000
w_sum_translation[1] = 000_10111100001111011100000
w_carry_translation[1] = 111_00110100010100000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01011110000111101110000 +
	110_10011010001010000000000
) = 2 * 111_11111000010001101110000 = 
111_11110000100011011100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_01111000011110111000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_01101000101000000000000
w_sum_translation[2] = 001_01111000011110111000000
w_carry_translation[2] = 110_01101000101000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	111_11110000100011011100000 +
	000_00000000000000000000000
) = 2 * 111_11110000100011011100000 = 
111_11100001000110111000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_11110000111101110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_11010001010000000000000
w_sum_translation[3] = 000_11110000111101110000000
w_carry_translation[3] = 110_11010001010000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	111_11100001000110111000000 +
	000_00000000000000000000000
) = 2 * 111_11100001000110111000000 = 
111_11000010001101110000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_11100001111011100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
101_10100010100000000000000
w_sum_translation[4] = 111_11100001111011100000000
w_carry_translation[4] = 111_10100010100000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_11 -> q[5] = -1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	111_11000010001101110000000 +
	000_00000000000000000000000
) = 2 * 111_11000010001101110000000 = 
111_10000100011011100000000
q_pos = 1000_0
q_neg = 0000_1

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
010_01001101011011000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_10000111001000000000000
w_sum_translation[5] = 000_01001101011011000000000
w_carry_translation[5] = 001_10000111001000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_01 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	111_10000100011011100000000 +
	001_01100101110110000000000
) = 2 * 000_11101010010001100000000 = 
001_11010100100011000000000
q_pos = 1000_01
q_neg = 0000_10


w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
110_10100000110010000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_00111100101000000000000
w_sum_translation[6] = 000_10100000110010000000000
w_carry_translation[6] = 000_00111100101000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 00_00 -> q[7] = +1
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	001_11010100100011000000000 +
	110_10011010001010000000000
) = 2 * 000_01101110101101000000000 = 
000_11011101011010000000000
q_pos = 1000_011
q_neg = 0000_100

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
100_00001100100000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_11100010101000000000000
w_sum_translation[7] = 110_00001100100000000000000
w_carry_translation[7] = 000_11100010101000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 10_00 -> q[8] = 0
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_11011101011010000000000 +
	110_10011010001010000000000
) = 2 * 111_01110111100100000000000 = 
110_11101111001000000000000
q_pos = 1000_0110
q_neg = 0000_1000

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	110_11101111001000000000000 +
	000_00000000000000000000000
) = 2 * 110_11101111001000000000000 = 
101_11011110010000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 000000111101001111111000 = 250872
D[WIDTH-1:0] = 000000000000000010111010 = 186
Q[WIDTH-1:0] = X / D = 1348 = 000000000000010101000100
REM[WIDTH-1:0] = 250872 - 186 * 1348 = 144 = 000000000000000010010000

CLZ_X = 6
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 10
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 12
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111101001111111000000000
Divisor[WIDTH-1:0] 		= 101110100000000000000000

+ D[(WIDTH + 2)-1:0] = 001_01110100000000000000000
+2D[(WIDTH + 2)-1:0] = 010_11101000000000000000000
- D[(WIDTH + 2)-1:0] = 110_10001100000000000000000
-2D[(WIDTH + 2)-1:0] = 101_00011000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[12];
w[final] = 110_10110000000000000000000 < 0
// 最后一次迭代的商
q[12] = 0
q_pos = 1011_0000_1100
q_neg = 0000_1000_0010
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
101010001010
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 10101000100
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1_10101100000000000000000 + 1_01110100000000000000000 = 
100100000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
100100000000000000000000 >> 16 = 
000000000000000010010000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_11101001111111000000000
w_sum_translation[0] = w_sum[0] =  001_01011110000111101110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

// 规格化之后必然有:
// q[1] = 1
// 为了方便人工计算，在草稿中一般可以直接令w_carry[1] = -2D, 实际的RTL实现中，是不知道-2D的值的(因为需要对D进行取反，然后再进行一个WIDTH宽度的全加操作).
w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_11010011111110000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_00011000000000000000000
w_sum_translation[1] = 001_11010011111110000000000
w_carry_translation[1] = 111_00011000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11101001111111000000000 +
	110_10001100000000000000000
) = 2 * 000_01110101111111000000000 = 
000_11101011111110000000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_10100111111100000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_00110000000000000000000
w_sum_translation[2] = 001_10100111111100000000000
w_carry_translation[2] = 000_00110000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_00 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_11101011111110000000000 +
	000_00000000000000000000000
) = 2 * 000_11101011111110000000000 = 
001_11010111111100000000000
q_pos = 101
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_00110111111000000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_10010000000000000000000
w_sum_translation[3] = 000_00110111111000000000000
w_carry_translation[3] = 000_10010000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_00 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_11010111111100000000000 +
	110_10001100000000000000000
) = 2 * 000_01100011111100000000000 = 
000_11000111111000000000000
q_pos = 1011
q_neg = 0000


w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_01010111110000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_01010000000000000000000
w_sum_translation[4] = 000_01010111110000000000000
w_carry_translation[4] = 110_01010000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_11000111111000000000000 +
	110_10001100000000000000000
) = 2 * 111_01010011111000000000000 = 
110_10100111110000000000000
q_pos = 1011_0
q_neg = 0000_0
abs(w[4]) = 001_01011000010000000000000
+D = 001_01110100000000000000000

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_10101111100000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_10100000000000000000000
w_sum_translation[5] = 110_10101111100000000000000
w_carry_translation[5] = 110_10100000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 10_10 -> q[6] = -2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	110_10100111110000000000000 +
	000_00000000000000000000000
) = 2 * 110_10100111110000000000000 = 
101_01001111100000000000000
q_pos = 1011_00
q_neg = 0000_10

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_11001111000000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_10100000000000000000000
w_sum_translation[6] = 111_11001111000000000000000
w_carry_translation[6] = 000_10100000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 11_00 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	101_01001111100000000000000 +
	010_11101000000000000000000
) = 2 * 000_00110111100000000000000 = 
000_01101111000000000000000
q_pos = 1011_000
q_neg = 0000_100

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_10011110000000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
001_01000000000000000000000
w_sum_translation[7] = 111_10011110000000000000000
w_carry_translation[7] = 001_01000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 11_01 -> q[8] = 0
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_01101111000000000000000 +
	000_00000000000000000000000
) = 2 * 000_01101111000000000000000 = 
000_11011110000000000000000
q_pos = 1011_0000
q_neg = 0000_1000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
111_00111100000000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
010_10000000000000000000000
w_sum_translation[8] = 001_00111100000000000000000
w_carry_translation[8] = 000_10000000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 01_00 -> q[9] = +1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	000_11011110000000000000000 +
	000_00000000000000000000000
) = 2 * 000_11011110000000000000000 = 
001_10111100000000000000000
q_pos = 1011_0000_1
q_neg = 0000_1000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
010_01100000000000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_00110000000000000000000
w_sum_translation[9] = 000_01100000000000000000000
w_carry_translation[9] = 000_00110000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_00 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	001_10111100000000000000000 +
	110_10001100000000000000000
) = 2 * 000_01001000000000000000000 = 
000_10010000000000000000000
q_pos = 1011_0000_11
q_neg = 0000_1000_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_10111000000000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
100_10000000000000000000000
w_sum_translation[10] = 111_10111000000000000000000
w_carry_translation[10] = 110_10000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 11_10 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	000_10010000000000000000000 +
	110_10001100000000000000000
) = 2 * 111_00011100000000000000000 = 
110_00111000000000000000000
q_pos = 1011_0000_110
q_neg = 0000_1000_001

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_10011000000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
010_11000000000000000000000
w_sum_translation[11] = 110_10011000000000000000000
w_carry_translation[11] = 000_11000000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_00 -> q[12] = 0
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	110_00111000000000000000000 +
	001_01110100000000000000000
) = 2 * 111_10101100000000000000000 = 
111_01011000000000000000000
q_pos = 1011_0000_1100
q_neg = 0000_1000_0010

// 最后一次迭代的余数
w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	111_01011000000000000000000 +
	000_00000000000000000000000
) = 2 * 111_01011000000000000000000 = 
110_10110000000000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 010110000000001111000111 = 5768135
D[WIDTH-1:0] = 000000100000000000000011 = 131075
Q[WIDTH-1:0] = X / D = 44 = 000000000000000000101100
REM[WIDTH-1:0] = 5768135 - 131075 * 44 = 835 = 000000000000001101000011

CLZ_X = 1
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 5
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 7
规格化操作之后:
Dividend[WIDTH-1:0] 	= 101100000000011110001110
Divisor[WIDTH-1:0] 		= 100000000000000011000000

+ D[(WIDTH + 2)-1:0] = 001_00000000000000011000000
+2D[(WIDTH + 2)-1:0] = 010_00000000000000110000000
- D[(WIDTH + 2)-1:0] = 110_11111111111111101000000
-2D[(WIDTH + 2)-1:0] = 101_11111111111111010000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[7];
w[final] = 000_00000110100001100000000 >= 0
// 最后一次迭代的商
q[7] = +2
q_pos = 1011_000
q_neg = 0000_000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
1011000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 101100
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
000000001101000011000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
000000001101000011000000 >> 6 = 
000000000000001101000011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 010110000000001111000111 = 5768135
D[WIDTH-1:0] = 000001000000000000000110 = 262150
Q[WIDTH-1:0] = X / D = 22 = 000000000000000000010110
REM[WIDTH-1:0] = 5768135 - 262150 * 22 = 835 = 000000000000001101000011

CLZ_X = 1
CLZ_D = 5
CLZ_DIFF = CLZ_D - CLZ_X = 4
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 6
w_sum_translation[5] = 000_00000001110110101000000
w_carry_translation[5] = 001_11111111110010100000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	010_00000000110100111100000 +
	110_11111111111111101000000
) = 2 * 001_00000000110100100100000 = 
010_00000001101001001000000
q_pos = 1011_00
q_neg = 0000_00
q_pos - q_neg = 00101100
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	010_00000001101001001000000 +
	101_11111111111111010000000
) = 2 * 000_00000001101000011000000 = 
000_00000011010000110000000

000_00000011010000110000000 / 4 = 000_00000000110100001100000
000000000110100001100000 >> CLZ_D = 000000000110100001100000 >> 5 =
000000000000001101000011
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_01100000000011110001110
w_sum_translation[0] = w_sum[0] =  001_01100000000011110001110
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0


w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_11000000000111100011100
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11111111111111010000000
w_sum_translation[1] = 000_11000000000111100011100
w_carry_translation[1] = 111_11111111111111010000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_01100000000011110001110 +
	110_11111111111111101000000
) = 2 * 000_01100000000011011001110 = 
000_11000000000110110011100
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_10000000001111000111000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11111111111110100000000
w_sum_translation[2] = 001_10000000001111000111000
w_carry_translation[2] = 111_11111111111110100000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_11000000000110110011100 +
	000_00000000000000000000000
) = 2 * 000_11000000000110110011100 = 
001_10000000001101100111000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_00000000011110001110000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_11111111111101000000000
w_sum_translation[3] = 001_00000000011110001110000
w_carry_translation[3] = 001_11111111111101000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_01 -> q[4] = +2
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_10000000001101100111000 +
	000_00000000000000000000000
) = 2 * 001_10000000001101100111000 = 
011_00000000011011001110000
q_pos = 1010
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_00000000111000111100000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11111111111100000000000
w_sum_translation[4] = 000_00000000111000111100000
w_carry_translation[4] = 001_11111111111100000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_01 -> q[5] = +1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	011_00000000011011001110000 +
	101_11111111111111010000000
) = 2 * 001_00000000011010011110000 = 
010_00000000110100111100000
q_pos = 1010_1
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_00000001110110101000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11111111110010100000000
w_sum_translation[5] = 000_00000001110110101000000
w_carry_translation[5] = 001_11111111110010100000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_01 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	010_00000000110100111100000 +
	110_11111111111111101000000
) = 2 * 001_00000000110100100100000 = 
010_00000001101001001000000
q_pos = 1010_11
q_neg = 0000_00


w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
110_00000011110111000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_11111111011010100000000
w_sum_translation[6] = 000_00000011110111000000000
w_carry_translation[6] = 001_11111111011010100000000
// 最后一次使用特殊的选择函数:
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 00_01 -> q[7] = +2
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	010_00000001101001001000000 +
	110_11111111111111101000000
) = 2 * 001_00000001101000110000000 = 
010_00000011010001100000000
q_pos = 1011_000
q_neg = 0000_000


w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	010_00000011010001100000000 +
	101_11111111111111010000000
) = 2 * 000_00000011010000110000000 = 
000_00000110100001100000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 001000000010011111110011 = 2107379
D[WIDTH-1:0] = 000000111111110000110000 = 261168
Q[WIDTH-1:0] = X / D = 8 = 000000000000000000001000
REM[WIDTH-1:0] = 2107379 - 261168 * 8 = 18035 = 000000000100011001110011

CLZ_X = 2
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 4
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 6
规格化操作之后:
Dividend[WIDTH-1:0] 	= 100000001001111111001100
Divisor[WIDTH-1:0] 		= 111111110000110000000000

+ D[(WIDTH + 2)-1:0] = 001_11111110000110000000000
+2D[(WIDTH + 2)-1:0] = 011_11111100001100000000000
- D[(WIDTH + 2)-1:0] = 110_00000001111010000000000
-2D[(WIDTH + 2)-1:0] = 100_00000011110100000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 000_10001100111001100000000 >= 0
// 最后一次迭代的商
q[6] = 0
q_pos = 1000_00
q_neg = 0100_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
00010000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0001000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
000100011001110011000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
000100011001110011000000 >> 6 = 
000000000100011001110011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 001000000010011111110011 = 2107379
D[WIDTH-1:0] = 001111111100001100000000 = 4178688
Q[WIDTH-1:0] = X / D = 0 = 000000000000000000000000
REM[WIDTH-1:0] = 2107379 - 4178688 * 0 = 2107379 = 001000000010011111110011

CLZ_X = 2
CLZ_D = 2
CLZ_DIFF = CLZ_D - CLZ_X = 0
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 2

// 最后一次迭代的余数
w[final] = w[2];
w[final] = 100_00001100100111100110000 < 0
// 最后一次迭代的商
q[2] = 0
q_pos = 10
q_neg = 00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
10
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1_00000011001001111001100 + 1_11111110000110000000000 = 
100000001001111111001100
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
100000001001111111001100 >> 2 = 
001000000010011111110011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 2)-1:0] =  001_00000001001111111001100
w_sum_translation[0] = w_sum[0] =  001_00000001001111111001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_00000010011111110011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_00000011110100000000000
w_sum_translation[1] = 000_00000010011111110011000
w_carry_translation[1] = 110_00000011110100000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_00000001001111111001100 +
	110_00000001111010000000000
) = 2 * 111_00000011001001111001100 = 
110_00000110010011110011000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_00000100111111100110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_00000111101000000000000
w_sum_translation[2] = 
w_carry_translation[2] = 
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 10_10 -> q[3] = -2
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_00000110010011110011000 +
	000_00000000000000000000000
) = 2 * 110_00000110010011110011000 = 
100_00001100100111100110000
q_pos = 100
q_neg = 010

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11111110110111001100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_00010010110000000000000
w_sum_translation[3] = 001_11111110110111001100000
w_carry_translation[3] = 110_00010010110000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	100_00001100100111100110000 +
	011_11111100001100000000000
) = 2 * 000_00001000110011100110000 = 
000_00010001100111001100000
q_pos = 1000
q_neg = 0100

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11111101101110011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_00100101100000000000000
w_sum_translation[4] = 001_11111101101110011000000
w_carry_translation[4] = 110_00100101100000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00010001100111001100000 +
	000_00000000000000000000000
) = 2 * 000_00010001100111001100000 = 
000_00100011001110011000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11111011011100110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_01001011000000000000000
w_sum_translation[5] = 001_11111011011100110000000
w_carry_translation[5] = 110_01001011000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_00100011001110011000000 +
	000_00000000000000000000000
) = 2 * 000_00100011001110011000000 = 
000_01000110011100110000000
q_pos = 1000_00
q_neg = 0100_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_11110110111001100000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
100_10010110000000000000000
w_sum_translation[6] = 001_11110110111001100000000
w_carry_translation[6] = 110_10010110000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_10 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_01000110011100110000000 +
	000_00000000000000000000000
) = 2 * 000_01000110011100110000000 = 
000_10001100111001100000000
q_pos = 1000_000
q_neg = 0100_000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 001111111111111110000011 = 4194179
D[WIDTH-1:0] = 000000000010000000110000 = 8240
Q[WIDTH-1:0] = X / D = 509 = 000000000000000111111101
REM[WIDTH-1:0] = 4194179 - 8240 * 509 = 19 = 000000000000000000010011

CLZ_X = 2
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 8
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 10
规格化操作之后:
Dividend[WIDTH-1:0] 	= 111111111111111000001100
Divisor[WIDTH-1:0] 		= 100000001100000000000000

+ D[(WIDTH + 2)-1:0] = 001_00000001100000000000000
+2D[(WIDTH + 2)-1:0] = 010_00000011000000000000000
- D[(WIDTH + 2)-1:0] = 110_11111110100000000000000
-2D[(WIDTH + 2)-1:0] = 101_11111101000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[10];
w[final] = 010_00000101011000000000000 >= 0
q[9] = +2
// 最后一次迭代的商
q[10] = +1
q_pos = 1111_1110_01
q_neg = 0000_0000_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 001111111001
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 111111100 -> 有问题, LSB比正确结果少1

出问题的原因在于(w[10] / 2)属于区间"[+D, +2D)"

// 先不管商的话, 如果使用另一种方法则能求出正确的余数
w[final] / 2 = 010_00000101011000000000000 / 2 = 100000010101100000000000
100000010101100000000000 + (-D) = 
100000010101100000000000 + 100000001100000000000000 = 
000000001001100000000000
000000001001100000000000 >> (CLZ_D + 1) = 000000001001100000000000 >> 11 = 000000000000000000010011

记住这一次的错误!!!!

// 出现了错误的结果...
// _??_
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
最后一次使用特殊的商选择函数, 使:
{w_sum_translation[i][MSB-1:MSB-2], w_carry_translation[i][MSB-1:MSB-2]} = 00_01, 01_00, 时选择q[i+1] = +2
{w_sum_translation[i][MSB-1:MSB-2], w_carry_translation[i][MSB-1:MSB-2]} = 11_10, 10_11, 时选择q[i+1] = -2
则有:
w_sum_translation[9] = 000_00110000001100000000000
w_carry_translation[9] = 001_11010100000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_01 -> q[10] = +2
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	011_00000101000110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000010000110000000000 = 
010_00000100001100000000000
q_pos = 1111_1110_10
q_neg = 0000_0000_00

w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	010_00000100001100000000000 +
	101_11111101000000000000000
) = 2 * 000_00000001001100000000000 = 
000_00000010011000000000000

// 最后一次迭代的余数
w[final] = w[10];
w[final] = 000_00000010011000000000000 >= 0
// 最后一次迭代的商
q_pos = 1111_1110_10
q_neg = 0000_0000_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
001111111010
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 00111111101
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
000000000100110000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
000000000100110000000000 >> 10 = 
000000000000000000010011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 001111111111111110000011 = 4194179
D[WIDTH-1:0] = 000001000000011000000000 = 263680
Q[WIDTH-1:0] = X / D = 15 = 000000000000000000001111
REM[WIDTH-1:0] = 4194179 - 263680 * 15 = 238979 = 000000111010010110000011

CLZ_X = 2
CLZ_D = 5
CLZ_DIFF = CLZ_D - CLZ_X = 3
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 5

w_sum_translation[4] = 001_11100001110000011000000
w_carry_translation[4] = 001_11110100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[5] = +2
q_pos = 1111_0
q_neg = 0000_0
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
11110
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[5] < 0))[WIDTH:1] = 1111

w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	011_11010101110000011000000 +
	101_11111101000000000000000
) = 2 * 001_11010010110000011000000 = 
011_10100101100000110000000

w[5] / 4 = 011_10100101100000110000000 / 4 = 011101001011000001100000
011101001011000001100000 >> CLZ_D = 011101001011000001100000 >> 5 = 
000000111010010110000011


// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 测试子集
X[WIDTH-1:0] = 001111111111111110000011 = 4194179
D[WIDTH-1:0] = 000000001000000011000000 = 32960
Q[WIDTH-1:0] = X / D = 127 = 000000000000000001111111
REM[WIDTH-1:0] = 4194179 - 32960 * 127 = 8259 = 000000000010000001000011

CLZ_X = 2
CLZ_D = 8
CLZ_DIFF = CLZ_D - CLZ_X = 6
多迭代一次, 迭代次数:
iter_num = CLZ_DIFF + 2 = 8

q[8] = +1
q_pos = 1111_1101
q_neg = 0000_0000
q_pos - q_neg = 11111101

w[8] = 011_00000101000110000000000 >= 0
w[8] / 2 = 001_10000010100011000000000
001_10000010100011000000000 + (-D) = 
001_10000010100011000000000 + 110_11111110100000000000000 = 
000_10000001000011000000000

010000001000011000000000 >> (CLZ_D + 1) = 
000000000010000001000011

// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 2)-1:0] =  001_11111111111111000001100
w_sum_translation[0] = w_sum[0] =  001_11111111111111000001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_11111111111110000011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11111101000000000000000
w_sum_translation[1] = 001_11111111111110000011000
w_carry_translation[1] = 111_11111101000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_11111111111111000001100 +
	110_11111110100000000000000
) = 2 * 000_11111110011111000001100 = 
001_11111100111110000011000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_11111111111100000110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_11111010000000000000000
w_sum_translation[2] = 001_11111111111100000110000
w_carry_translation[2] = 001_11111010000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_01 -> q[3] = +2
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	001_11111100111110000011000 +
	000_00000000000000000000000
) = 2 * 001_11111100111110000011000 = 
011_11111001111100000110000
q_pos = 110
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_11110001111000001100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11111100000000000000000
w_sum_translation[3] = 001_11110001111000001100000
w_carry_translation[3] = 001_11111100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_01 -> q[4] = +2
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	011_11111001111100000110000 +
	101_11111101000000000000000
) = 2 * 001_11110110111100000110000 = 
011_11101101111000001100000
q_pos = 1110
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_11100001110000011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11110100000000000000000
w_sum_translation[4] = 001_11100001110000011000000
w_carry_translation[4] = 001_11110100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_01 -> q[5] = +2
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	011_11101101111000001100000 +
	101_11111101000000000000000
) = 2 * 001_11101010111000001100000 = 
011_11010101110000011000000
q_pos = 1111_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_11010001100000110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_11010100000000000000000
w_sum_translation[5] = 001_11010001100000110000000
w_carry_translation[5] = 001_11010100000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	011_11010101110000011000000 +
	101_11111101000000000000000
) = 2 * 001_11010010110000011000000 = 
011_10100101100000110000000
q_pos = 1111_10
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_11110001000001100000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_01010100000000000000000
w_sum_translation[6] = 001_11110001000001100000000
w_carry_translation[6] = 001_01010100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_01 -> q[7] = +2
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_10100101100000110000000 +
	101_11111101000000000000000
) = 2 * 001_10100010100000110000000 = 
011_01000101000001100000000
q_pos = 1111_110
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_10110000000011000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
011_11010100000000000000000
w_sum_translation[7] = 000_10110000000011000000000
w_carry_translation[7] = 001_11010100000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	011_01000101000001100000000 +
	101_11111101000000000000000
) = 2 * 001_01000010000001100000000 = 
010_10000100000011000000000
q_pos = 1111_1101
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
111_00110101000110000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
011_11010000000000000000000
w_sum_translation[8] = 001_00110101000110000000000
w_carry_translation[8] = 001_11010000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 01_01 -> q[9] = +2
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	010_10000100000011000000000 +
	110_11111110100000000000000
) = 2 * 001_10000010100011000000000 = 
011_00000101000110000000000
q_pos = 1111_1110_0
q_neg = 0000_0000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_00110000001100000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
011_11010100000000000000000
w_sum_translation[9] = 000_00110000001100000000000
w_carry_translation[9] = 001_11010100000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 00_01 -> q[10] = +1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	011_00000101000110000000000 +
	101_11111101000000000000000
) = 2 * 001_00000010000110000000000 = 
010_00000100001100000000000
q_pos = 1111_1110_01
q_neg = 0000_0000_00


w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
110_00110101011000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
011_11010000000000000000000
w_sum_translation[10] = 000_00110101011000000000000
w_carry_translation[10] = 001_11010000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 00_01 -> q[11] = +1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	010_00000100001100000000000 +
	110_11111110100000000000000
) = 2 * 001_00000010101100000000000 = 
010_00000101011000000000000
q_pos = 1111_1110_011
q_neg = 0000_0000_000

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
110_00110111110000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
011_11010000000000000000000
w_sum_translation[11] = 000_00110111110000000000000
w_carry_translation[11] = 001_11010000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 00_01 -> q[12] = +1
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	010_00000101011000000000000 +
	110_11111110100000000000000
) = 2 * 001_00000011111000000000000 = 
010_00000111110000000000000
q_pos = 1111_1110_0111
q_neg = 0000_0000_0000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 001000000110011111110011 = 2123763
D[WIDTH-1:0] = 000000111111110000000001 = 261121
Q[WIDTH-1:0] = X / D = 8 = 000000000000000000001000
REM[WIDTH-1:0] = 2123763 - 261121 * 8 = 34795 = 000000001000011111101011

CLZ_X = 2
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 4
迭代次数:
iter_num = CLZ_DIFF + 1 + 1 = 6
规格化操作之后:
Dividend[WIDTH-1:0] 	= 100000011001111111001100
Divisor[WIDTH-1:0] 		= 111111110000000001000000

+ D[(WIDTH + 2)-1:0] = 001_11111110000000001000000
+2D[(WIDTH + 2)-1:0] = 011_11111100000000010000000
- D[(WIDTH + 2)-1:0] = 110_00000001111111111000000
-2D[(WIDTH + 2)-1:0] = 100_00000011111111110000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 001_00001111110101100000000 >= 0
// 最后一次迭代的商
q[6] = 0
q_pos = 1000_00
q_neg = 0100_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
00010000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0001000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[WIDTH-1:0] + (w[final] < 0 ? D[WIDTH-1:0] : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
0_01000011111101011000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
001000011111101011000000 >> 6 = 
000000001000011111101011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 2)-1:0] =  001_00000011001111111001100
w_sum_translation[0] = w_sum[0] =  001_00000011001111111001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_00000000000000000000000
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_00000110011111110011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_00000011111111110000000
w_sum_translation[1] = 000_00000110011111110011000
w_carry_translation[1] = 110_00000011111111110000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_00000011001111111001100 +
	110_00000001111111111000000
) = 2 * 111_00000101001111110001100 = 
110_00001010011111100011000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_00001100111111100110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_00000111111111100000000
w_sum_translation[2] = 110_00001100111111100110000
w_carry_translation[2] = 110_00000111111111100000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 10_10 -> q[3] = -2
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_00001010011111100011000 +
	000_00000000000000000000000
) = 2 * 110_00001010011111100011000 = 
100_00010100111111000110000
q_pos = 100
q_neg = 010

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11101110000000101100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_00110011111110000000000
w_sum_translation[3] = 001_11101110000000101100000
w_carry_translation[3] = 110_00110011111110000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	100_00010100111111000110000 +
	011_11111100000000010000000
) = 2 * 000_00010000111111010110000 = 
000_00100001111110101100000
q_pos = 1000
q_neg = 0100

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_11011100000001011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_01100111111100000000000
w_sum_translation[4] = 001_11011100000001011000000
w_carry_translation[4] = 110_01100111111100000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00100001111110101100000 +
	000_00000000000000000000000
) = 2 * 000_00100001111110101100000 = 
000_01000011111101011000000
q_pos = 1000_0
q_neg = 0100_0


w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_10111000000010110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_11001111111000000000000
w_sum_translation[5] = 001_10111000000010110000000
w_carry_translation[5] = 110_11001111111000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_01000011111101011000000 +
	000_00000000000000000000000
) = 2 * 000_01000011111101011000000 = 
000_10000111111010110000000
q_pos = 1000_00
q_neg = 0100_00

w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_10000111111010110000000 +
	000_00000000000000000000000
) = 2 * 000_10000111111010110000000 = 
001_00001111110101100000000







// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 32;
ITN = InTerNal
ITN_W = 1 + WIDTH = 33;
0_00000000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 10000001010111000000011000101110 = 2170291758
D[WIDTH-1:0] = 00000001001101000001100110100011 = 20191651
Q[WIDTH-1:0] = X / D = 107 = 00000000000000000000000001101011
REM[WIDTH-1:0] = 2170291758 - 20191651 * 107 = 9785101 = 00000000100101010100111100001101

CLZ_X = 0
CLZ_D = 7
CLZ_DIFF = CLZ_D - CLZ_X = 7
Normalized_D = 10011010000011001101000110000000
根据D的值, 可得选择常数:
m[-1] = -14
m[ 0] = - 4
m[+1] = + 4
m[+2] = +14

+ D[ITN_W-1:0] = 0_10011010000011001101000110000000
+2D[ITN_W-1:0] = 1_00110100000110011010001100000000
- D[ITN_W-1:0] = 1_01100101111100110010111010000000
-2D[ITN_W-1:0] = 0_11001011111001100101110100000000
~ D[ITN_W-1:0] = 1_01100101111100110010111001111111
~2D[ITN_W-1:0] = 0_11001011111001100101110011111111

l_shift_num = CLZ_D = 7
shifted_dividend[(2 * WIDTH + 1)-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_0000000000000000000000000000000010000001010111000000011000101110 << 7 = 
0_0000000000000000000000000100000010101110000000110001011100000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w_sum[0][ITN_W-1:0] 	= 0_00000000000000000000000001000000
w_carry[0][ITN_W-1:0] 	= 0_00000000000000000000000000000000
w[0] 					= 0_00000000000000000000000001000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
10101110000000110001011100000000

ITER[0]:
w_sum[1] = csa_sum({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000100000010
w_carry[1] = csa_carry({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000000000000
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_00000000000000000000000100000010 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000000100000010
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
10111000000011000101110000000000

ITER[1]:
w_sum[2] = csa_sum({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000010000001010
w_carry[2] = csa_carry({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000000000000000
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_00000000000000000000010000001010 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000010000001010
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
11100000001100010111000000000000

ITER[2]:
w_sum[3] = csa_sum({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000001000000101011
w_carry[3] = csa_carry({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000000000000000
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_00000000000000000001000000101011 + 
0_00000000000000000000000000000000 = 
0_00000000000000000001000000101011
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
10000000110001011100000000000000

ITER[3]:
w_sum[4] = csa_sum({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000100000010101110
w_carry[4] = csa_carry({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000000000000000000
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_00000000000000000100000010101110 + 
0_00000000000000000000000000000000 = 
0_00000000000000000100000010101110
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
00000011000101110000000000000000

ITER[4]:
w_sum[5] = csa_sum({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000010000001010111000
w_carry[5] = csa_carry({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000000000000000000000
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_00000000000000010000001010111000 + 
0_00000000000000000000000000000000 = 
0_00000000000000010000001010111000
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
00001100010111000000000000000000

ITER[5]:
w_sum[6] = csa_sum({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000001000000101011100000
w_carry[6] = csa_carry({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000000000000000000000000
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_00000000000001000000101011100000 + 
0_00000000000000000000000000000000 = 
0_00000000000001000000101011100000
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
00110001011100000000000000000000

ITER[6]:
w_sum[7] = csa_sum({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000100000010101110000000
w_carry[7] = csa_carry({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000000000000000000000000
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_00000000000100000010101110000000 + 
0_00000000000000000000000000000000 = 
0_00000000000100000010101110000000
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
11000101110000000000000000000000

ITER[7]:
w_sum[8] = csa_sum({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000010000001010111000000011
w_carry[8] = csa_carry({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000000000000000000000000000
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_00000000010000001010111000000011 + 
0_00000000000000000000000000000000 = 
0_00000000010000001010111000000011
(4 * w[8])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
(4 * w_sum[8])_trunc_3_4 + (4 * w_carry[8])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
00010111000000000000000000000000

ITER[8]:
w_sum[9] = csa_sum({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000001000000101011100000001100
w_carry[9] = csa_carry({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000000000000000000000000000000
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_00000001000000101011100000001100 + 
0_00000000000000000000000000000000 = 
0_00000001000000101011100000001100
(4 * w[9])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
(4 * w_sum[9])_trunc_3_4 + (4 * w_carry[9])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
01011100000000000000000000000000

ITER[9]:
w_sum[10] = csa_sum({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000100000010101110000000110001
w_carry[10] = csa_carry({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000000000000000000000000000000
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_00000100000010101110000000110001 + 
0_00000000000000000000000000000000 = 
0_00000100000010101110000000110001
(4 * w[10])_trunc_3_4 = 000_0001, "belongs to [m[0], m[+1])" -> q[11] = 0
(4 * w_sum[10])_trunc_3_4 + (4 * w_carry[10])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[0], m[+1])" -> q[11] = 0
q_pos = 0000_0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
01110000000000000000000000000000

ITER[10]:
w_sum[11] = csa_sum({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00010000001010111000000011000101
w_carry[11] = csa_carry({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00000000000000000000000000000000
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
0_00010000001010111000000011000101 + 
0_00000000000000000000000000000000 = 
0_00010000001010111000000011000101
(4 * w[11])_trunc_3_4 = 000_0100, "belongs to [m[+1], m[+2])" -> q[12] = +1
(4 * w_sum[11])_trunc_3_4 + (4 * w_carry[11])_trunc_3_4 = 
000_0100 + 000_0000 = 000_0100, "belongs to [m[+1], m[+2])" -> q[12] = +1
q_pos = 0000_0000_0000_0000_0000_0001
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
11000000000000000000000000000000

ITER[11]:
w_sum[12] = csa_sum({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
1_00100101010111010010110101101000
w_carry[12] = csa_carry({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
0_10000001010001000000010000101111
w[12] = {w[11] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[12] * D = 
0_01000000101011100000001100010111 + 
1_01100101111100110010111010000000 = 
1_10100110101000010011000110010111
(4 * w[12])_trunc_3_4 = 110_1001, "belongs to [-Inf, m[-1])" -> q[13] = -2
(4 * w_sum[12])_trunc_3_4 + (4 * w_carry[12])_trunc_3_4 = 
100_1001 + 010_0000 = 110_1001, "belongs to [-Inf, m[-1])" -> q[13] = -2
q_pos = 0000_0000_0000_0000_0000_0001_00
q_neg = 0000_0000_0000_0000_0000_0000_10
temp_dividend[12] = temp_dividend[11] << 2 = 
00000000000000000000000000000000
\
ITER[12]:
w_sum[13] = csa_sum({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
1_10100100011111010000011000011100
w_carry[13] = csa_carry({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
0_00101010001000010110001101000000
w[13] = {w[12] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[13] * D = 
0_10011010100001001100011001011100 + 
1_00110100000110011010001100000000 = 
1_11001110100111100110100101011100
(4 * w[13])_trunc_3_4 = 111_0011, "belongs to [m[-1], m[0])" -> q[14] = -1
(4 * w_sum[13])_trunc_3_4 + (4 * w_carry[13])_trunc_3_4 = 
110_1001 + 000_1010 = 111_0011, "belongs to [m[-1], m[0])" -> q[14] = -1
q_pos = 0000_0000_0000_0000_0000_0001_0000
q_neg = 0000_0000_0000_0000_0000_0000_1001
temp_dividend[13] = temp_dividend[12] << 2 = 
00000000000000000000000000000000

ITER[13]:
w_sum[14] = csa_sum({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
0_10100011011111010100010011110000
w_carry[14] = csa_carry({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
1_00110001000010010011001000000000
w[14] = {w[13] << 2, temp_dividend[12][(WIDTH-1) -: 2]} - q[14] * D = 
1_00111010011110011010010101110000 + 
0_10011010000011001101000110000000 = 
1_11010100100001100111011011110000
(4 * w[14])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[15] = -1
(4 * w_sum[14])_trunc_3_4 + (4 * w_carry[14])_trunc_3_4 = 
010_1000 + 100_1100 = 111_0100, "belongs to [m[-1], m[0])" -> q[15] = -1
q_pos = 0000_0000_0000_0000_0000_0001_0000_00
q_neg = 0000_0000_0000_0000_0000_0000_1001_01
temp_dividend[14] = temp_dividend[13] << 2 = 
00000000000000000000000000000000

ITER[14]:
w_sum[15] = csa_sum({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
0_11010011110111010000101001000000
w_carry[15] = csa_carry({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
1_00011000010010011010001100000000
w[15] = {w[14] << 2, temp_dividend[13][(WIDTH-1) -: 2]} - q[15] * D = 
1_01010010000110011101101111000000 + 
0_10011010000011001101000110000000 = 
1_11101100001001101010110101000000
(4 * w[15])_trunc_3_4 = 111_1011, "belongs to [m[-1], m[0])" -> q[16] = -1
(4 * w_sum[15])_trunc_3_4 + (4 * w_carry[15])_trunc_3_4 = 
011_0100 + 100_0110 = 111_1010, "belongs to [m[-1], m[0])" -> q[16] = -1
q_pos = 0000_0000_0000_0000_0000_0001_0000_0000
q_neg = 0000_0000_0000_0000_0000_0000_1001_0101
temp_dividend[15] = temp_dividend[14] << 2 = 
00000000000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w_sum[16] = csa_sum({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
1_10110100010111100111010010000000
w_carry[16] = csa_carry({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
0_10010110010010010001001000000000
w[16] = {w[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]} - q[16] * D = 
1_10110000100110101011010100000000 + 
0_10011010000011001101000110000000 = 
0_01001010101001111000011010000000 >= 0



rem = (w[final])_trunc >> CLZ_D = 
01001010101001111000011010000000 >> 7 = 
00000000100101010100111100001101

q_final = corr(q_pos - q_neg) = 01101011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 01010101100001100101010100010101 = 1434866965
D[WIDTH-1:0] = 00000010000101100011100110010010 = 35010962
Q[WIDTH-1:0] = X / D = 40 = 00000000000000000000000000101000
REM[WIDTH-1:0] = 1434866965 - 35010962 * 40 = 34428485 = 00000010000011010101011001000101

CLZ_X = 0
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 6
Normalized_D = 10000101100011100110010010000000
根据D的值, 可得选择常数:
m[-1] = -14
m[ 0] = - 4
m[+1] = + 4
m[+2] = +14

+ D[ITN_W-1:0] = 0_10000101100011100110010010000000
+2D[ITN_W-1:0] = 1_00001011000111001100100100000000
- D[ITN_W-1:0] = 1_01111010011100011001101110000000
-2D[ITN_W-1:0] = 0_11110100111000110011011100000000
~ D[ITN_W-1:0] = 1_01111010011100011001101101111111
~2D[ITN_W-1:0] = 0_11110100111000110011011011111111

l_shift_num = CLZ_D = 6
shifted_dividend[(2 * WIDTH + 1)-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_0000000000000000000000000000000001010101100001100101010100010101 << 6 = 
0_0000000000000000000000000001010101100001100101010100010101000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w_sum[0][ITN_W-1:0] 	= 0_00000000000000000000000000010101
w_carry[0][ITN_W-1:0] 	= 0_00000000000000000000000000000000
w[0] 					= 0_00000000000000000000000000010101
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
01100001100101010100010101000000

ITER[0]:
w_sum[1] = csa_sum({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000001010101
w_carry[1] = csa_carry({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000000000000
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_00000000000000000000000001010101 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000000001010101
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
10000110010101010001010100000000

ITER[1]:
w_sum[2] = csa_sum({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000000101010110
w_carry[2] = csa_carry({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000000000000000
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_00000000000000000000000101010110 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000000101010110
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
00011001010101000101010000000000

ITER[2]:
w_sum[3] = csa_sum({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000010101011000
w_carry[3] = csa_carry({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000000000000000
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_00000000000000000000010101011000 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000010101011000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
01100101010100010101000000000000

ITER[3]:
w_sum[4] = csa_sum({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000001010101100001
w_carry[4] = csa_carry({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000000000000000000
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_00000000000000000001010101100001 + 
0_00000000000000000000000000000000 = 
0_00000000000000000001010101100001
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
10010101010001010100000000000000

ITER[4]:
w_sum[5] = csa_sum({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000000101010110000110
w_carry[5] = csa_carry({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000000000000000000000
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_00000000000000000101010110000110 + 
0_00000000000000000000000000000000 = 
0_00000000000000000101010110000110
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
01010101000101010000000000000000

ITER[5]:
w_sum[6] = csa_sum({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000000010101011000011001
w_carry[6] = csa_carry({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000000000000000000000000
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_00000000000000010101011000011001 + 
0_00000000000000000000000000000000 = 
0_00000000000000010101011000011001
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
01010100010101000000000000000000

ITER[6]:
w_sum[7] = csa_sum({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000001010101100001100101
w_carry[7] = csa_carry({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000000000000000000000000
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_00000000000001010101100001100101 + 
0_00000000000000000000000000000000 = 
0_00000000000001010101100001100101
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
01010001010100000000000000000000

ITER[7]:
w_sum[8] = csa_sum({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000000101010110000110010101
w_carry[8] = csa_carry({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000000000000000000000000000
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_00000000000101010110000110010101 + 
0_00000000000000000000000000000000 = 
0_00000000000101010110000110010101
(4 * w[8])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
(4 * w_sum[8])_trunc_3_4 + (4 * w_carry[8])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
01000101010000000000000000000000

ITER[8]:
w_sum[9] = csa_sum({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000000010101011000011001010101
w_carry[9] = csa_carry({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000000000000000000000000000000
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_00000000010101011000011001010101 + 
0_00000000000000000000000000000000 = 
0_00000000010101011000011001010101
(4 * w[9])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
(4 * w_sum[9])_trunc_3_4 + (4 * w_carry[9])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
00010101000000000000000000000000

ITER[9]:
w_sum[10] = csa_sum({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000001010101100001100101010100
w_carry[10] = csa_carry({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000000000000000000000000000000
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_00000001010101100001100101010100 + 
0_00000000000000000000000000000000 = 
0_00000001010101100001100101010100
(4 * w[10])_trunc_3_4 = 000_0001, "belongs to [m[0], m[+1])" -> q[11] = 0
(4 * w_sum[10])_trunc_3_4 + (4 * w_carry[10])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[0], m[+1])" -> q[11] = 0
q_pos = 0000_0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
01010100000000000000000000000000

ITER[10]:
w_sum[11] = csa_sum({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00000101010110000110010101010001
w_carry[11] = csa_carry({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00000000000000000000000000000000
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
0_00000101010110000110010101010001 + 
0_00000000000000000000000000000000 = 
0_00000101010110000110010101010001
(4 * w[11])_trunc_3_4 = 000_0001, "belongs to [m[+1], m[+2])" -> q[12] = 0
(4 * w_sum[11])_trunc_3_4 + (4 * w_carry[11])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[+1], m[+2])" -> q[12] = 0
q_pos = 0000_0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
01010000000000000000000000000000

ITER[11]:
w_sum[12] = csa_sum({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
0_00010101011000011001010101000101
w_carry[12] = csa_carry({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
0_00000000000000000000000000000000
w[12] = {w[11] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[12] * D = 
0_00010101011000011001010101000101 + 
0_00000000000000000000000000000000 = 
0_00010101011000011001010101000101
(4 * w[12])_trunc_3_4 = 000_0101, "belongs to [m[+1], m[+2])" -> q[13] = +1
(4 * w_sum[12])_trunc_3_4 + (4 * w_carry[12])_trunc_3_4 = 
000_0101 + 000_0000 = 000_0101, "belongs to [m[+1], m[+2])" -> q[13] = +1
q_pos = 0000_0000_0000_0000_0000_0000_01
q_neg = 0000_0000_0000_0000_0000_0000_00
temp_dividend[12] = temp_dividend[11] << 2 = 
01000000000000000000000000000000

ITER[12]:
w_sum[13] = csa_sum({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
1_00101111111101111100111001101010
w_carry[13] = csa_carry({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
0_10100000000000000010001000101011
w[13] = {w[12] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[13] * D = 
0_01010101100001100101010100010101 + 
1_01111010011100011001101110000000 = 
1_11001111111101111111000010010101
(4 * w[13])_trunc_3_4 = 111_0011, "belongs to [m[-1], m[0])" -> q[14] = -1
(4 * w_sum[13])_trunc_3_4 + (4 * w_carry[13])_trunc_3_4 = 
100_1011 + 010_1000 = 111_0011, "belongs to [m[-1], m[0])" -> q[14] = -1
q_pos = 0000_0000_0000_0000_0000_0000_0100
q_neg = 0000_0000_0000_0000_0000_0000_0001
temp_dividend[13] = temp_dividend[12] << 2 = 
00000000000000000000000000000000

ITER[13]:
w_sum[14] = csa_sum({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
0_10111010010100011101010110000100
w_carry[14] = csa_carry({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
1_00001011000111000101000101010000
w[14] = {w[13] << 2, temp_dividend[12][(WIDTH-1) -: 2]} - q[14] * D = 
1_00111111110111111100001001010100 + 
0_10000101100011100110010010000000 = 
1_11000101011011100010011011010100
(4 * w[14])_trunc_3_4 = 111_0001, "belongs to [-Inf, m[-1])" -> q[15] = -2
(4 * w_sum[14])_trunc_3_4 + (4 * w_carry[14])_trunc_3_4 = 
010_1110 + 100_0010 = 111_0000, "belongs to [-Inf, m[-1])" -> q[15] = -2
q_pos = 0000_0000_0000_0000_0000_0000_0100_00
q_neg = 0000_0000_0000_0000_0000_0000_0001_10
temp_dividend[14] = temp_dividend[13] << 2 = 
00000000000000000000000000000000

ITER[14]:
w_sum[15] = csa_sum({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
1_11001110001010101101101001010000
w_carry[15] = csa_carry({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
0_01010010101010101000101000000000
w[15] = {w[14] << 2, temp_dividend[13][(WIDTH-1) -: 2]} - q[15] * D = 
1_00010101101110001001101101010000 + 
1_00001011000111001100100100000000 = 
0_00100000110101010110010001010000
(4 * w[15])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[16] = +1
(4 * w_sum[15])_trunc_3_4 + (4 * w_carry[15])_trunc_3_4 = 
111_0011 + 001_0100 = 000_0111, "belongs to [m[+1], m[+2])" -> q[16] = +1
q_pos = 0000_0000_0000_0000_0000_0000_0100_0001
q_neg = 0000_0000_0000_0000_0000_0000_0001_1000
temp_dividend[15] = temp_dividend[14] << 2 = 
00000000000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w_sum[16] = csa_sum({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
1_00001000011100001101101000111111
w_carry[16] = csa_carry({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
0_11110101010101100101001010000001
w[16] = {w[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]} - q[16] * D = 
0_10000011010101011001000101000000 + 
1_01111010011100011001101110000000 = 
1_11111101110001110010110011000000 < 0


rem = (w[final] + D)_trunc >> CLZ_D = 
(11111101110001110010110011000000 + 10000101100011100110010010000000) >> 6 = 
10000011010101011001000101000000 >> 6 = 
00000010000011010101011001000101

q_final = corr(q_pos - q_neg) = 00101000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 10100011010010000010001000100001 = 2739413537
D[WIDTH-1:0] = 00000010111110010100111101100010 = 49893218
Q[WIDTH-1:0] = X / D = 54 = 00000000000000000000000000110110
REM[WIDTH-1:0] = 2739413537 - 49893218 * 54 = 45179765 = 00000010101100010110001101110101

CLZ_X = 0
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 6
Normalized_D = 10111110010100111101100010000000
根据D的值, 可得选择常数:
m[-1] = -16
m[ 0] = - 6
m[+1] = + 6
m[+2] = +16

+ D[ITN_W-1:0] = 0_10111110010100111101100010000000
+2D[ITN_W-1:0] = 1_01111100101001111011000100000000
- D[ITN_W-1:0] = 1_01000001101011000010011110000000
-2D[ITN_W-1:0] = 0_10000011010110000100111100000000
~ D[ITN_W-1:0] = 1_01000001101011000010011101111111
~2D[ITN_W-1:0] = 0_10000011010110000100111011111111

l_shift_num = CLZ_D = 6
shifted_dividend[(2 * WIDTH + 1)-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_0000000000000000000000000000000010100011010010000010001000100001 << 6 = 
0_0000000000000000000000000010100011010010000010001000100001000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w_sum[0][ITN_W-1:0] 	= 0_00000000000000000000000000101000
w_carry[0][ITN_W-1:0] 	= 0_00000000000000000000000000000000
w[0] 					= 0_00000000000000000000000000101000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00
temp_dividend[0][WIDTH-1:0] = shifted_dividend[WIDTH-1:0] = 
11010010000010001000100001000000

ITER[0]:
w_sum[1] = csa_sum({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000010100011
w_carry[1] = csa_carry({w_sum[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]}, 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000000000000
w[1] = {w[0] << 2, temp_dividend[0][(WIDTH-1) -: 2]} - q[1] * D = 
0_00000000000000000000000010100011 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000000010100011
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000
temp_dividend[1] = temp_dividend[0] << 2 = 
01001000001000100010000100000000

ITER[1]:
w_sum[2] = csa_sum({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000001010001101
w_carry[2] = csa_carry({w_sum[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]}, 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000000000000000
w[2] = {w[1] << 2, temp_dividend[1][(WIDTH-1) -: 2]} - q[2] * D = 
0_00000000000000000000001010001101 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000001010001101
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00
temp_dividend[2] = temp_dividend[1] << 2 = 
00100000100010001000010000000000

ITER[2]:
w_sum[3] = csa_sum({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000101000110100
w_carry[3] = csa_carry({w_sum[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]}, 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000000000000000
w[3] = {w[2] << 2, temp_dividend[2][(WIDTH-1) -: 2]} - q[3] * D = 
0_00000000000000000000101000110100 + 
0_00000000000000000000000000000000 = 
0_00000000000000000000101000110100
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000
temp_dividend[3] = temp_dividend[2] << 2 = 
10000010001000100001000000000000

ITER[3]:
w_sum[4] = csa_sum({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000010100011010010
w_carry[4] = csa_carry({w_sum[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]}, 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000000000000000000
w[4] = {w[3] << 2, temp_dividend[3][(WIDTH-1) -: 2]} - q[4] * D = 
0_00000000000000000010100011010010 + 
0_00000000000000000000000000000000 = 
0_00000000000000000010100011010010
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00
temp_dividend[4] = temp_dividend[3] << 2 = 
00001000100010000100000000000000

ITER[4]:
w_sum[5] = csa_sum({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000001010001101001000
w_carry[5] = csa_carry({w_sum[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]}, 4 * w_carry[4], -q[5] * D) = 
0_00000000000000000000000000000000
w[5] = {w[4] << 2, temp_dividend[4][(WIDTH-1) -: 2]} - q[5] * D = 
0_00000000000000001010001101001000 + 
0_00000000000000000000000000000000 = 
0_00000000000000001010001101001000
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000
temp_dividend[5] = temp_dividend[4] << 2 = 
00100010001000010000000000000000

ITER[5]:
w_sum[6] = csa_sum({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000000101000110100100000
w_carry[6] = csa_carry({w_sum[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]}, 4 * w_carry[5], -q[6] * D) = 
0_00000000000000000000000000000000
w[6] = {w[5] << 2, temp_dividend[5][(WIDTH-1) -: 2]} - q[6] * D = 
0_00000000000000101000110100100000 + 
0_00000000000000000000000000000000 = 
0_00000000000000101000110100100000
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00
temp_dividend[6] = temp_dividend[5] << 2 = 
10001000100001000000000000000000

ITER[6]:
w_sum[7] = csa_sum({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000010100011010010000010
w_carry[7] = csa_carry({w_sum[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]}, 4 * w_carry[6], -q[7] * D) = 
0_00000000000000000000000000000000
w[7] = {w[6] << 2, temp_dividend[6][(WIDTH-1) -: 2]} - q[7] * D = 
0_00000000000010100011010010000010 + 
0_00000000000000000000000000000000 = 
0_00000000000010100011010010000010
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000
temp_dividend[7] = temp_dividend[6] << 2 = 
00100010000100000000000000000000

ITER[7]:
w_sum[8] = csa_sum({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000001010001101001000001000
w_carry[8] = csa_carry({w_sum[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]}, 4 * w_carry[7], -q[8] * D) = 
0_00000000000000000000000000000000
w[8] = {w[7] << 2, temp_dividend[7][(WIDTH-1) -: 2]} - q[8] * D = 
0_00000000001010001101001000001000 + 
0_00000000000000000000000000000000 = 
0_00000000001010001101001000001000
(4 * w[8])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
(4 * w_sum[8])_trunc_3_4 + (4 * w_carry[8])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00
temp_dividend[8] = temp_dividend[7] << 2 = 
10001000010000000000000000000000

ITER[8]:
w_sum[9] = csa_sum({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000000101000110100100000100010
w_carry[9] = csa_carry({w_sum[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]}, 4 * w_carry[8], -q[9] * D) = 
0_00000000000000000000000000000000
w[9] = {w[8] << 2, temp_dividend[8][(WIDTH-1) -: 2]} - q[9] * D = 
0_00000000101000110100100000100010 + 
0_00000000000000000000000000000000 = 
0_00000000101000110100100000100010
(4 * w[9])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
(4 * w_sum[9])_trunc_3_4 + (4 * w_carry[9])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[10] = 0
q_pos = 0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000
temp_dividend[9] = temp_dividend[8] << 2 = 
00100001000000000000000000000000

ITER[9]:
w_sum[10] = csa_sum({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000010100011010010000010001000
w_carry[10] = csa_carry({w_sum[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]}, 4 * w_carry[9], -q[10] * D) = 
0_00000000000000000000000000000000
w[10] = {w[9] << 2, temp_dividend[9][(WIDTH-1) -: 2]} - q[10] * D = 
0_00000010100011010010000010001000 + 
0_00000000000000000000000000000000 = 
0_00000010100011010010000010001000
(4 * w[10])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[11] = 0
(4 * w_sum[10])_trunc_3_4 + (4 * w_carry[10])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[0], m[+1])" -> q[11] = 0
q_pos = 0000_0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_0000_00
temp_dividend[10] = temp_dividend[9] << 2 = 
10000100000000000000000000000000

ITER[10]:
w_sum[11] = csa_sum({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00001010001101001000001000100010
w_carry[11] = csa_carry({w_sum[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]}, 4 * w_carry[10], -q[11] * D) = 
0_00000000000000000000000000000000
w[11] = {w[10] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[11] * D = 
0_00001010001101001000001000100010 + 
0_00000000000000000000000000000000 = 
0_00001010001101001000001000100010
(4 * w[11])_trunc_3_4 = 000_0010, "belongs to [m[+1], m[+2])" -> q[12] = 0
(4 * w_sum[11])_trunc_3_4 + (4 * w_carry[11])_trunc_3_4 = 
000_0010 + 000_0000 = 000_0010, "belongs to [m[+1], m[+2])" -> q[12] = 0
q_pos = 0000_0000_0000_0000_0000_0000
q_neg = 0000_0000_0000_0000_0000_0000
temp_dividend[11] = temp_dividend[10] << 2 = 
00010000000000000000000000000000

ITER[11]:
w_sum[12] = csa_sum({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
0_00101000110100100000100010001000
w_carry[12] = csa_carry({w_sum[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]}, 4 * w_carry[11], -q[12] * D) = 
0_00000000000000000000000000000000
w[12] = {w[11] << 2, temp_dividend[10][(WIDTH-1) -: 2]} - q[12] * D = 
0_00101000110100100000100010001000 + 
0_00000000000000000000000000000000 = 
0_00101000110100100000100010001000
(4 * w[12])_trunc_3_4 = 000_1010, "belongs to [m[+1], m[+2])" -> q[13] = +1
(4 * w_sum[12])_trunc_3_4 + (4 * w_carry[12])_trunc_3_4 = 
000_1010 + 000_0000 = 000_1010, "belongs to [m[+1], m[+2])" -> q[13] = +1
q_pos = 0000_0000_0000_0000_0000_0000_01
q_neg = 0000_0000_0000_0000_0000_0000_00
temp_dividend[12] = temp_dividend[11] << 2 = 
01000000000000000000000000000000

ITER[12]:
w_sum[13] = csa_sum({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
1_11100010111001000000010101011110
w_carry[13] = csa_carry({w_sum[12] << 2, temp_dividend[12][(WIDTH-1) -: 2]}, 4 * w_carry[12], -q[13] * D) = 
0_00000010000100000100010001000011
w[13] = {w[12] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[13] * D = 
0_10100011010010000010001000100001 + 
1_01000001101011000010011110000000 = 
1_11100100111101000100100110100001
(4 * w[13])_trunc_3_4 = 111_1001, "belongs to [m[-1], m[0])" -> q[14] = -1
(4 * w_sum[13])_trunc_3_4 + (4 * w_carry[13])_trunc_3_4 = 
111_1000 + 000_0000 = 111_1000, "belongs to [m[-1], m[0])" -> q[14] = -1
q_pos = 0000_0000_0000_0000_0000_0000_0100
q_neg = 0000_0000_0000_0000_0000_0000_0001
temp_dividend[13] = temp_dividend[12] << 2 = 
00000000000000000000000000000000

ITER[13]:
w_sum[14] = csa_sum({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
1_00111101100000101101110011110100
w_carry[14] = csa_carry({w_sum[13] << 2, temp_dividend[13][(WIDTH-1) -: 2]}, 4 * w_carry[13], -q[14] * D) = 
1_00010100101000100010001000010000
w[14] = {w[13] << 2, temp_dividend[12][(WIDTH-1) -: 2]} - q[14] * D = 
1_10010011110100010010011010000100 + 
0_10111110010100111101100010000000 = 
0_01010010001001001111111100000100
(4 * w[14])_trunc_3_4 = 001_0100, "belongs to [m[+2], +Inf)" -> q[15] = +2
(4 * w_sum[14])_trunc_3_4 + (4 * w_carry[14])_trunc_3_4 = 
100_1111 + 100_0101 = 001_0100, "belongs to [m[+2], +Inf)" -> q[15] = +2
q_pos = 0000_0000_0000_0000_0000_0000_0100_10
q_neg = 0000_0000_0000_0000_0000_0000_0001_00
temp_dividend[14] = temp_dividend[13] << 2 = 
00000000000000000000000000000000

ITER[14]:
w_sum[15] = csa_sum({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
0_00100111110110111011010101101111
w_carry[15] = csa_carry({w_sum[14] << 2, temp_dividend[14][(WIDTH-1) -: 2]}, 4 * w_carry[14], -q[15] * D) = 
1_10100100000100001001010110100001
w[15] = {w[14] << 2, temp_dividend[13][(WIDTH-1) -: 2]} - q[15] * D = 
1_01001000100100111111110000010000 + 
0_10000011010110000100111100000000 = 
1_11001011111011000100101100010000
(4 * w[15])_trunc_3_4 = 111_0010, "belongs to [m[-1], m[0])" -> q[16] = -1
(4 * w_sum[15])_trunc_3_4 + (4 * w_carry[15])_trunc_3_4 = 
000_1001 + 110_1001 = 111_0010, "belongs to [m[-1], m[0])" -> q[16] = -1
q_pos = 0000_0000_0000_0000_0000_0000_0100_1000
q_neg = 0000_0000_0000_0000_0000_0000_0001_0001
temp_dividend[15] = temp_dividend[14] << 2 = 
00000000000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w_sum[16] = csa_sum({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
0_10110001011111110101101110111000
w_carry[16] = csa_carry({w_sum[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]}, 4 * w_carry[15], -q[16] * D) = 
1_00111100100001011010100100001000
w[16] = {w[15] << 2, temp_dividend[15][(WIDTH-1) -: 2]} - q[16] * D = 
1_00101111101100010010110001000000 + 
0_10111110010100111101100010000000 = 
1_11101110000001010000010011000000 < 0


rem = (w[final] + D)_trunc >> CLZ_D = 
(11101110000001010000010011000000 + 10111110010100111101100010000000) >> 6 = 
10101100010110001101110101000000 >> 6 = 
00000010101100010110001101110101

q_final = corr(q_pos - q_neg) = 00110110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


















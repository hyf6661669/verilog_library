测试不移位的Non-Restoring除法, 在操作数位宽较小的时候此算法可能会有优势。



// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 24
// ---------------------------------------------------------------------------------------------------------------------------------------
// TODO
X[WIDTH-1:0] = 000010101111000011110111 = 717047
D[WIDTH-1:0] = 000000000000000010101011 = 171
Q[WIDTH-1:0] = X / D = 4193 = 000000000001000001100001
REM[WIDTH-1:0] = 717047 - 171 * 4193 = 44 = 000000000000000000101100

CLZ_X = 4
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 12
迭代次数:
iter_num = CLZ_DIFF + 1 = 13

+D = 101010110000000000000000

初始化:
rem[0] 	= 101011110000111101110000
d[0] 	= 101010110000000000000000
q[0] = 0

ITER[0]:
rem[1] = rem[0] + (q[0] ? -d[0] : d[0]) = 
101011110000111101110000 + 
-101010110000000000000000 = 
000001000000111101110000 >= 0 -> q[1] = 1

d[1] = d[0] >> 1 = 010101011000000000000000
rem[2] = rem[1] + (q[1] ? -d[1] : d[1]) = 
000001000000111101110000 + 
-010101011000000000000000 = 
101011101000111101110000 < 0 -> q[2] = 0

d[2] = d[1] >> 1 = 001010101100000000000000
rem[3] = rem[2] + (q[2] ? -d[2] : d[2]) = 
101011101000111101110000 + 
001010101100000000000000 = 
110110010100111101110000 < 0 -> q[3] = 0

d[3] = d[2] >> 1 = 000101010110000000000000
rem[4] = rem[3] + (q[3] ? -d[3] : d[3]) = 
110110010100111101110000 + 
000101010110000000000000 = 
111011101010111101110000 < 0 -> q[4] = 0

d[4] = d[3] >> 1 = 000010101011000000000000
rem[5] = rem[4] + (q[4] ? -d[4] : d[4]) = 
111011101010111101110000 + 
000010101011000000000000 = 
111110010101111101110000 < 0 -> q[5] = 0

d[5] = d[4] >> 1 = 000001010101100000000000
rem[6] = rem[5] + (q[5] ? -d[5] : d[5]) = 
111110010101111101110000 + 
000001010101100000000000 = 
111111101011011101110000 < 0 -> q[6] = 0

d[6] = d[5] >> 1 = 000000101010110000000000
rem[7] = rem[6] + (q[6] ? -d[6] : d[6]) = 
111111101011011101110000 + 
000000101010110000000000 = 
000000010110001101110000 >= 0 -> q[7] = 1

d[7] = d[6] >> 1 = 000000010101011000000000
rem[8] = rem[7] + (q[7] ? -d[7] : d[7]) = 
000000010110001101110000 + 
-000000010101011000000000 = 
000000000000110101110000 >= 0 -> q[8] = 1

d[8] = d[7] >> 1 = 000000001010101100000000
rem[9] = rem[8] + (q[8] ? -d[8] : d[8]) = 
000000000000110101110000 + 
-000000001010101100000000 = 
111111110110001001110000 < 0 -> q[9] = 0

d[9] = d[8] >> 1 = 000000000101010110000000
rem[10] = rem[9] + (q[9] ? -d[9] : d[9]) = 
111111110110001001110000 + 
000000000101010110000000 = 
111111111011011111110000 < 0 -> q[10] = 0

d[10] = d[9] >> 1 = 000000000010101011000000
rem[11] = rem[10] + (q[10] ? -d[10] : d[10]) = 
111111111011011111110000 + 
000000000010101011000000 = 
111111111110001010110000 < 0 -> q[11] = 0

d[11] = d[10] >> 1 = 000000000001010101100000
rem[12] = rem[11] + (q[11] ? -d[11] : d[11]) = 
111111111110001010110000 + 
000000000001010101100000 = 
111111111111100000010000 < 0 -> q[12] = 0

d[12] = d[11] >> 1 = 000000000000101010110000
rem[13] = rem[12] + (q[12] ? -d[12] : d[12]) = 
111111111111100000010000 + 
000000000000101010110000 = 
000000000000001011000000 >= 0 -> q[13] = 1


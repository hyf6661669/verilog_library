!!!!!!注意!!!!!!
下面的例子里右移的方法似乎有误, 详见别的文档.


接"test_broken_0.sv", 此处探究的内容:
将1个或多个"Over-Redundant Radix-2"串联起来形成"High-Radix"除法器时，应该如何操作才能得到正确的余数.
对于Radix-N来说, 将Dividend变换到区间"[1, 2)"上之后, 需要再向右移:
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N));
N =  4 -> r_shift_num = 1 - ((CLZ_DIFF + 1) % 2);
N =  8 -> r_shift_num = 2 - ((CLZ_DIFF + 1) % 3);
N = 16 -> r_shift_num = 3 - ((CLZ_DIFF + 1) % 4);
N = 32 -> r_shift_num = 4 - ((CLZ_DIFF + 1) % 5);
N = 64 -> r_shift_num = 6 - ((CLZ_DIFF + 1) % 6);

这样最后一次"Radix-N"迭代计算出的"(log2(N))-bit"的商刚好是Q[0 +: log2(N)].
按照上述方法, 做WIDTH-bit整数除法时, 需要用(WIDTH + 2 + log2(N) - 1) = (WIDTH + 1 + log2(N))来表示w[i].
WIDTH = 28;

// ---------------------------------------------------------------------------------------------------------------------------------------
注意!!!!!!
在这个文件里的例子中发现了一个求余数时的注意事项，如果最后一次迭代为:
q[final] = -1/+1;
则应当使用如下方法计算remainder:
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 2)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0];
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> (CLZ_D + 1) = 
即不再是除以4, 而是应该除以2了.
自己分析的原因:
q[final] = -1/+1时, 说明最后一次的商应当比实际选中的商还要小1, 即:
q_correct[final] = q[final] - 1 -> q_correct[final] = -2/0;
所以将余数由负数恢复到正数时, 就需要将"w[final] / 2", 然后再加上"Divisor"来得到正的余数。
另一种情况里:
q[final] = -2/0/+2;
则说明"q_calculated_pre[0] = 0", 所以"q_calculated_pre - 1'b1"会将"q_calculated_pre[1]"减去1, 那么这个"- 1'b1"的操作等价于说明, 为了得到正的余数
需要把q[final - 1]减去1, 那么此时就需要将"w[final] / 4", 然后再加上"Divisor"来得到正的余数。
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
将3个Radix-2串联起来形成Radix-8算法, 即:
N = 8;
(WIDTH + 1 + log2(N)) = 32;

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110100001110011100100011 = 13690659
D[WIDTH-1:0] = 0000000000010010011101110111 = 75639
Q[WIDTH-1:0] = X / D = 181 = 0000000000000000000010110101
REM[WIDTH-1:0] = 13690659 - 75639 * 181 = 0 = 0000000000000000000000000000

CLZ_X = 4
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 7
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 2 - (8 % 3) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(9 / 3) = 3;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1101000011100111001000110000
Divisor[WIDTH-1:0] 		= 1001001110111011100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00100111011101110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_01001110111011100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11011000100010010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_10110001000100100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[9];
w[final] = 000_00000000000000000000000000000 >= 0
// 最后一次迭代的商
q[9] = 0
q_pos = 1011_0101_0
q_neg = 0000_0000_0
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
101101010
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 10110101
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
0000000000000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0000000000000000000000000000 >> 11 = 
0000000000000000000000000000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_10100001110011100100011000000
w_sum_translation[0] = w_sum[0] =  001_10100001110011100100011000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_01000011100111001000110000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_10110001000100100000000000000
w_sum_translation[1] = 001_01000011100111001000110000000
w_carry_translation[1] = 111_10110001000100100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_10100001110011100100011000000 +
	110_11011000100010010000000000000
) = 2 * 000_01111010010101110100011000000 = 
000_11110100101011101000110000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
010_10000111001110010001100000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_01100010001001000000000000000
w_sum_translation[2] = 000_10000111001110010001100000000
w_carry_translation[2] = 001_01100010001001000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_01 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_11110100101011101000110000000 +
	000_00000000000000000000000000000
) = 2 * 000_11110100101011101000110000000 = 
001_11101001010111010001100000000
q_pos = 101
q_neg = 000

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_01111011001010000011000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_00001000101001000000000000000
w_sum_translation[3] = 000_01111011001010000011000000000
w_carry_translation[3] = 001_00001000101001000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_01 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_11101001010111010001100000000 +
	110_11011000100010010000000000000
) = 2 * 000_11000001111001100001100000000 = 
001_10000011110011000011000000000
q_pos = 1011
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_01010110000010100110000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_01100010101000000000000000000
w_sum_translation[4] = 111_01010110000010100110000000000
w_carry_translation[4] = 001_01100010101000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_01 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	001_10000011110011000011000000000 +
	110_11011000100010010000000000000
) = 2 * 000_01011100010101010011000000000 = 
000_10111000101010100110000000000
q_pos = 1011_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_10101100000101001100000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
010_11000101010000000000000000000
w_sum_translation[5] = 000_10101100000101001100000000000
w_carry_translation[5] = 000_11000101010000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_00 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_10111000101010100110000000000 +
	000_00000000000000000000000000000
) = 2 * 000_10111000101010100110000000000 = 
001_01110001010101001100000000000
q_pos = 1011_01
q_neg = 0000_00

// 第3次大迭代
w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_01100011101110111000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_00110000000000000000000000000
w_sum_translation[6] = 111_01100011101110111000000000000
w_carry_translation[6] = 001_00110000000000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 11_01 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	001_01110001010101001100000000000 +
	110_11011000100010010000000000000
) = 2 * 000_01001001110111011100000000000 = 
000_10010011101110111000000000000
q_pos = 1011_010
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_11000111011101110000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_01100000000000000000000000000
w_sum_translation[7] = 000_11000111011101110000000000000
w_carry_translation[7] = 000_01100000000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_00 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_10010011101110111000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_10010011101110111000000000000 = 
001_00100111011101110000000000000
q_pos = 1011_0101
q_neg = 0000_0000

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
100_11111111111111000000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
011_00000000000001000000000000000
w_sum_translation[8] = 110_11111111111111000000000000000
w_carry_translation[8] = 001_00000000000001000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_01 -> q[9] = 0
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	001_00100111011101110000000000000 +
	110_11011000100010010000000000000
) = 2 * 000_00000000000000000000000000000 = 
000_00000000000000000000000000000
q_pos = 1011_0101_0
q_neg = 0000_0000_0

w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	000_00000000000000000000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_00000000000000000000000000000 = 
000_00000000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000000010100010100001100001 = 665697
D[WIDTH-1:0] = 0000000000010011100001111111 = 79999
Q[WIDTH-1:0] = X / D = 8 = 0000000000000000000000001000
REM[WIDTH-1:0] = 665697 - 79999 * 8 = 25705 = 0000000000000110010001101001

CLZ_X = 8
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 3
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 2 - (4 % 3) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(5 / 3) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1010001010000110000100000000
Divisor[WIDTH-1:0] 		= 1001110000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00111000011111110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_01110000111111100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11000111100000010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_10001111000000100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 001_10010001101001000000000000000 >= 0
// 最后一次迭代的商
q[6] = 0
q_pos = 1000_00
q_neg = 0100_00
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
00010000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0001000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
110010001101001000000000000000 / 4 = 
001100100011010010000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0011001000110100100000000000 >> 11 = 
0000000000000110010001101001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_10100010100001100001000000000
w_sum_translation[0] = w_sum[0] =  000_10100010100001100001000000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
001_01000101000011000010000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_10001111000000100000000000000
w_sum_translation[1] = 111_01000101000011000010000000000
w_carry_translation[1] = 111_10001111000000100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_10100010100001100001000000000 +
	110_11000111100000010000000000000
) = 2 * 111_01101010000001110001000000000 = 
110_11010100000011100010000000000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_11100100111000100100000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_00110100001110000000000000000
w_sum_translation[2] = 001_11100100111000100100000000000
w_carry_translation[2] = 110_00110100001110000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_11010100000011100010000000000 +
	001_00111000011111110000000000000
) = 2 * 000_00001100100011010010000000000 = 
000_00011001000110100100000000000
q_pos = 100
q_neg = 010

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11001001110001001000000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_01101000011100000000000000000
w_sum_translation[3] = 001_11001001110001001000000000000
w_carry_translation[3] = 110_01101000011100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00011001000110100100000000000 +
	000_00000000000000000000000000000
) = 2 * 000_00011001000110100100000000000 = 
000_00110010001101001000000000000
q_pos = 1000
q_neg = 0100

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_10010011100010010000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_11010000111000000000000000000
w_sum_translation[4] = 001_10010011100010010000000000000
w_carry_translation[4] = 110_11010000111000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00110010001101001000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_00110010001101001000000000000 = 
000_01100100011010010000000000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_00100111000100100000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
101_10100001110000000000000000000
w_sum_translation[5] = 001_00100111000100100000000000000
w_carry_translation[5] = 111_10100001110000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_11 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_01100100011010010000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_01100100011010010000000000000 = 
000_11001000110100100000000000000
q_pos = 1000_00
q_neg = 0100_00

w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_11001000110100100000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_11001000110100100000000000000 = 
001_10010001101001000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000001000001011111100000010 = 2146050
D[WIDTH-1:0] = 0000000000010000100001111111 = 67711
Q[WIDTH-1:0] = X / D = 31 = 0000000000000000000000011111
REM[WIDTH-1:0] = 2146050 - 67711 * 31 = 47009 = 0000000000001011011110100001

CLZ_X = 6
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 5
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 2 - (6 % 3) = 2;
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(7 / 3) = 3;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000001011111100000010000000
Divisor[WIDTH-1:0] 		= 1000010000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00001000011111110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_00010000111111100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11110111100000010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_11101111000000100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[9];
w[final] = 110_10111100100010000000000000000 < 0
// 最后一次迭代的商
q[9] = -2
q_pos = 1000_0000_0
q_neg = 0110_0000_0
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
01000000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0011111
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1101011110010001000000000000 + 1000010000111111100000000000 = 
0101101111010000100000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0101101111010000100000000000 >> 11 = 
0000000000001011011110100001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_01000001011111100000010000000
w_sum_translation[0] = w_sum[0] =  000_01000001011111100000010000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_10000010111111000000100000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11101111000000100000000000000
w_sum_translation[1] = 110_10000010111111000000100000000
w_carry_translation[1] = 111_11101111000000100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_01000001011111100000010000000 +
	110_11110111100000010000000000000
) = 2 * 111_00111000111111110000010000000 = 
110_01110001111111100000100000000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_11001011000000100001000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_00101001111110000000000000000
w_sum_translation[2] = 000_11001011000000100001000000000
w_carry_translation[2] = 110_00101001111110000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_01110001111111100000100000000 +
	001_00001000011111110000000000000
) = 2 * 111_01111010011111010000100000000 = 
110_11110100111110100001000000000
q_pos = 100
q_neg = 010

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
001_10010110000001000010000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_01010011111100000000000000000
w_sum_translation[3] = 111_10010110000001000010000000000
w_carry_translation[3] = 110_01010011111100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_10 -> q[4] = -1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	110_11110100111110100001000000000 +
	000_00000000000000000000000000000
) = 2 * 110_11110100111110100001000000000 = 
101_11101001111101000010000000000
q_pos = 1000
q_neg = 0101

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_10011011000101100100000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_01001001110100000000000000000
w_sum_translation[4] = 111_10011011000101100100000000000
w_carry_translation[4] = 110_01001001110100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_10 -> q[5] = -1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	101_11101001111101000010000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11110010011100110010000000000 = 
101_11100100111001100100000000000
q_pos = 1000_0
q_neg = 0101_1

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
001_10110101011100101000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_00100101010110000000000000000
w_sum_translation[5] = 111_10110101011100101000000000000
w_carry_translation[5] = 110_00100101010110000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 11_10 -> q[6] = -1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	101_11100100111001100100000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11101101011001010100000000000 = 
101_11011010110010101000000000000
q_pos = 1000_00
q_neg = 0101_11

// 第3次大迭代
w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_00110000101010110000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
100_10010101111010000000000000000
w_sum_translation[6] = 111_00110000101010110000000000000
w_carry_translation[6] = 110_10010101111010000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 11_10 -> q[7] = -1
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	101_11011010110010101000000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11100011010010011000000000000 = 
101_11000110100100110000000000000
q_pos = 1000_000
q_neg = 0101_111

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
001_01011010011110000000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
100_01000011101011000000000000000
w_sum_translation[7] = 111_01011010011110000000000000000
w_carry_translation[7] = 110_01000011101011000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 11_10 -> q[8] = -1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	101_11000110100100110000000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11001111000100100000000000000 = 
101_10011110001001000000000000000
q_pos = 1000_0000
q_neg = 0101_1111

w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
000_00100011010101100000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
101_00101001111100000000000000000
w_sum_translation[8] = 110_00100011010101100000000000000
w_carry_translation[8] = 111_00101001111100000000000000000
// 最后一次迭代使用特殊的选择函数
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_11 -> q[9] = -2
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	101_10011110001001000000000000000 +
	001_00001000011111110000000000000
) = 2 * 110_10100110101000110000000000000 = 
101_01001101010001100000000000000
q_pos = 1000_0000_0
q_neg = 0110_0000_0

w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	101_01001101010001100000000000000 +
	010_00010000111111100000000000000
) = 2 * 111_01011110010001000000000000000 = 
110_10111100100010000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
将4个Radix-2串联起来形成Radix-16算法, 即:
N = 16;
(WIDTH + 1 + log2(N)) = 33;

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000010001100010111011110011 = 4599539
D[WIDTH-1:0] = 0000000000000001000111010100 = 4564
Q[WIDTH-1:0] = X / D = 1007 = 0000000000000000001111101111
REM[WIDTH-1:0] = 4599539 - 4564 * 1007 = 3591 = 0000000000000000111000000111

CLZ_X = 5
CLZ_D = 15
CLZ_DIFF = CLZ_D - CLZ_X = 10
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (11 % 4) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(12 / 4) = 3;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000110001011101111001100000
Divisor[WIDTH-1:0] 		= 1000111010100000000000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_000111010100000000000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_001110101000000000000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_111000101100000000000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_110001011000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[12];
w[final] = 111_000011001100000000000000000000 < 0
// 最后一次迭代的商
q[12] = -2
q_pos = 1000_0000_0000
q_neg = 0000_0010_0000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 
011111100000
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 01111101111
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1110000110011000000000000000 + 1000111010100000000000000000 = 
0111000000111000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0111000000111000000000000000 >> 15 = 
0000000000000000111000000111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_000110001011101111001100000000
w_sum_translation[0] = w_sum[0] =  001_000110001011101111001100000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_001100010111011110011000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_110001011000000000000000000000
w_sum_translation[1] = 000_001100010111011110011000000000
w_carry_translation[1] = 111_110001011000000000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_000110001011101111001100000000 +
	110_111000101100000000000000000000
) = 2 * 111_111110110111101111001100000000 = 
111_111101101111011110011000000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_011000101110111100110000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_100010110000000000000000000000
w_sum_translation[2] = 000_011000101110111100110000000000
w_carry_translation[2] = 111_100010110000000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	111_111101101111011110011000000000 +
	000_000000000000000000000000000000
) = 2 * 111_111101101111011110011000000000 = 
111_111011011110111100110000000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_110001011101111001100000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_000101100000000000000000000000
w_sum_translation[3] = 000_110001011101111001100000000000
w_carry_translation[3] = 111_000101100000000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	111_111011011110111100110000000000 +
	000_000000000000000000000000000000
) = 2 * 111_111011011110111100110000000000 = 
111_110110111101111001100000000000
q_pos = 1000
q_neg = 0000

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_100010111011110011000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_001011000000000000000000000000
w_sum_translation[4] = 001_100010111011110011000000000000
w_carry_translation[4] = 110_001011000000000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	111_110110111101111001100000000000 +
	000_000000000000000000000000000000
) = 2 * 111_110110111101111001100000000000 = 
111_101101111011110011000000000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_000101110111100110000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_010110000000000000000000000000
w_sum_translation[5] = 001_000101110111100110000000000000
w_carry_translation[5] = 110_010110000000000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	111_101101111011110011000000000000 +
	000_000000000000000000000000000000
) = 2 * 111_101101111011110011000000000000 = 
111_011011110111100110000000000000
q_pos = 1000_00
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_001011101111001100000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
100_101100000000000000000000000000
w_sum_translation[6] = 000_001011101111001100000000000000
w_carry_translation[6] = 110_101100000000000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 00_10 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	111_011011110111100110000000000000 +
	000_000000000000000000000000000000
) = 2 * 111_011011110111100110000000000000 = 
110_110111101111001100000000000000
q_pos = 1000_000
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
000_010111011110011000000000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
101_011000000000000000000000000000
w_sum_translation[7] = 110_010111011110011000000000000000
w_carry_translation[7] = 111_011000000000000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 10_11 -> q[8] = -1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	110_110111101111001100000000000000 +
	000_000000000000000000000000000000
) = 2 * 110_110111101111001100000000000000 = 
101_101111011110011000000000000000
q_pos = 1000_0000
q_neg = 0000_0001

// 第3次大迭代
w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
000_010000010100110000000000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
101_011101010000000000000000000000
w_sum_translation[8] = 110_010000010100110000000000000000
w_carry_translation[8] = 111_011101010000000000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_11 -> q[9] = -1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	101_101111011110011000000000000000 +
	001_000111010100000000000000000000
) = 2 * 110_110110110010011000000000000000 = 
101_101101100100110000000000000000
q_pos = 1000_0000_0
q_neg = 0000_0001_1

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
000_010100100001100000000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
101_010101010000000000000000000000
w_sum_translation[9] = 110_010100100001100000000000000000
w_carry_translation[9] = 111_010101010000000000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_11 -> q[10] = -1
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	101_101101100100110000000000000000 +
	001_000111010100000000000000000000
) = 2 * 110_110100111000110000000000000000 = 
101_101001110001100000000000000000
q_pos = 1000_0000_00
q_neg = 0000_0001_11

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
000_001101001011000000000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
101_010101000000000000000000000000
w_sum_translation[10] = 110_001101001011000000000000000000
w_carry_translation[10] = 111_010101000000000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 10_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	101_101001110001100000000000000000 +
	001_000111010100000000000000000000
) = 2 * 110_110001000101100000000000000000 = 
101_100010001011000000000000000000
q_pos = 1000_0000_000
q_neg = 0000_0001_111

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
000_111110111110000000000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
100_010100000000000000000000000000
w_sum_translation[11] = 110_111110111110000000000000000000
w_carry_translation[11] = 110_010100000000000000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 10_10 -> q[12] = -2
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	101_100010001011000000000000000000 +
	001_000111010100000000000000000000
) = 2 * 110_101001011111000000000000000000 = 
101_010010111110000000000000000000
q_pos = 1000_0000_0000
q_neg = 0000_0010_0000

w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	101_010010111110000000000000000000 +
	010_001110101000000000000000000000
) = 2 * 111_100001100110000000000000000000 = 
111_000011001100000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0111111111100010111011110011 = 134098675
D[WIDTH-1:0] = 0000001111110001000101000011 = 4133187
Q[WIDTH-1:0] = X / D = 32 = 0000000000000000000000100000
REM[WIDTH-1:0] = 134098675 - 4133187 * 32 = 1836691 = 0000000111000000011010010011

CLZ_X = 1
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 5
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (6 % 4) = 1;
迭代次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(7 / 4) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111111111000101110111100110
Divisor[WIDTH-1:0] 		= 1111110001000101000011000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_111110001000101000011000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 011_111100010001010000110000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_000001110111010111101000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 100_000011101110101111010000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8];
w[final] = 111_100011111011111000110000000000 < 0
// 最后一次迭代的商
q[7] = 0
q[final] = q[8] = +1
q_pos = 1000_0001
q_neg = 0100_0000
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 01000001
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0100000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 2)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1110001111101111100011000000 + 1111110001000101000011000000 = 
1110000000110100100110000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> (CLZ_D + 1) = 
1110000000110100100110000000 >> 7 = 
0000000111000000011010010011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_111111111100010111011110011000
w_sum_translation[0] = w_sum[0] =  000_111111111100010111011110011000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
001_111111111000101110111100110000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_000011101110101111010000000000
w_sum_translation[1] = 111_111111111000101110111100110000
w_carry_translation[1] = 110_000011101110101111010000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_10 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_111111111100010111011110011000 +
	110_000001110111010111101000000000
) = 2 * 111_000001110011101111000110011000 = 
110_000011100111011110001100110000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_000100111101010011101001100000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_111110100010111001100000000000
w_sum_translation[2] = 000_000100111101010011101001100000
w_carry_translation[2] = 111_111110100010111001100000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_000011100111011110001100110000 +
	001_111110001000101000011000000000
) = 2 * 000_000001110000000110100100110000 = 
000_000011100000001101001001100000
q_pos = 100
q_neg = 010

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_001001111010100111010011000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_111101000101110011000000000000
w_sum_translation[3] = 000_001001111010100111010011000000
w_carry_translation[3] = 111_111101000101110011000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_000011100000001101001001100000 +
	000_000000000000000000000000000000
) = 2 * 000_000011100000001101001001100000 = 
000_000111000000011010010011000000
q_pos = 1000
q_neg = 0100

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_010011110101001110100110000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_111010001011100110000000000000
w_sum_translation[4] = 000_010011110101001110100110000000
w_carry_translation[4] = 111_111010001011100110000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_11 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_000111000000011010010011000000 +
	000_000000000000000000000000000000
) = 2 * 000_000111000000011010010011000000 = 
000_001110000000110100100110000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_100111101010011101001100000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_110100010111001100000000000000
w_sum_translation[5] = 000_100111101010011101001100000000
w_carry_translation[5] = 111_110100010111001100000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_11 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_001110000000110100100110000000 +
	000_000000000000000000000000000000
) = 2 * 000_001110000000110100100110000000 = 
000_011100000001101001001100000000
q_pos = 1000_00
q_neg = 0100_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_001111010100111010011000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_101000101110011000000000000000
w_sum_translation[6] = 001_001111010100111010011000000000
w_carry_translation[6] = 111_101000101110011000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_11 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_011100000001101001001100000000 +
	000_000000000000000000000000000000
) = 2 * 000_011100000001101001001100000000 = 
000_111000000011010010011000000000
q_pos = 1000_000
q_neg = 0100_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_011110101001110100110000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_010001011100110000000000000000
w_sum_translation[7] = 000_011110101001110100110000000000
w_carry_translation[7] = 001_010001011100110000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_111000000011010010011000000000 +
	000_000000000000000000000000000000
) = 2 * 000_111000000011010010011000000000 = 
001_110000000110100100110000000000
q_pos = 1000_0001
q_neg = 0100_0000

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	001_110000000110100100110000000000 +
	110_000001110111010111101000000000
) = 2 * 111_110001111101111100011000000000 =
111_100011111011111000110000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0111111111100010111011110011 = 134098675
D[WIDTH-1:0] = 0000010000110001000101000011 = 4395331
Q[WIDTH-1:0] = X / D = 30 = 0000000000000000000000011110
REM[WIDTH-1:0] = 134098675 - 4395331 * 30 = 2238745 = 0000001000100010100100011001

CLZ_X = 1
CLZ_D = 5
CLZ_DIFF = CLZ_D - CLZ_X = 4
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (5 % 4) = 2;
迭代次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(6 / 4) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111111111000101110111100110
Divisor[WIDTH-1:0] 		= 1000011000100010100001100000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_000011000100010100001100000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_000110001000101000011000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_111100111011101011110100000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_111001110111010111101000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// TODO
// 最后一次迭代的余数
w[final] = w[8];
w[final] = 000_000010100000011101111000000000 >= 0
// 最后一次迭代的商
q[7] = 0
q[final] = q[8] = +1
q_pos = 1000_0001
q_neg = 0100_0100
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 00111101
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0011110
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 2)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
0000001010000001110111100000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> (CLZ_D + 1) = 
0000001010000001110111100000 >> 6 = 
0000000000001010000001110111
// _??_
又出错了!!!!

如果q[8] = 0:
q_pos = 1000_0000
q_neg = 0100_0100
q_calculated_pre = 00111100
q_calculated = 0011110
w[8] = 010_001000101001000110010000000000
w[8] / 4 = 0100010001010010001100100000
0100010001010010001100100000 >> 5 = 0000001000100010100100011001
这tmd倒是对了??
// _??_


000_000010100000011101111000000000 / 2 = 000_000001010000001110111100000000

000_000001010000001110111100000000 + D = 
000_000001010000001110111100000000 + 001_000011000100010100001100000000 = 
001_000100010100100011001000000000

001_000100010100100011001000000000 >> (CLZ_D + 1) = 
1000100010100100011001000000 >> 6 = 
0000001000100010100100011001


// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_011111111110001011101111001100
w_sum_translation[0] = w_sum[0] =  000_011111111110001011101111001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_111111111100010111011110011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_111001110111010111101000000000
w_sum_translation[1] = 110_111111111100010111011110011000
w_carry_translation[1] = 111_111001110111010111101000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_011111111110001011101111001100 +
	110_111100111011101011110100000000
) = 2 * 111_011100111001110111100011001100 = 
110_111001110011101111000110011000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_001010011110101001110100110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_101111010001011100110000000000
w_sum_translation[2] = 000_001010011110101001110100110000
w_carry_translation[2] = 111_101111010001011100110000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_111001110011101111000110011000 +
	001_000011000100010100001100000000
) = 2 * 111_111100111000000011010010011000 = 
111_111001110000000110100100110000
q_pos = 100
q_neg = 010

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_010100111101010011101001100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_011110100010111001100000000000
w_sum_translation[3] = 000_010100111101010011101001100000
w_carry_translation[3] = 111_011110100010111001100000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	111_111001110000000110100100110000 +
	000_000000000000000000000000000000
) = 2 * 111_111001110000000110100100110000 = 
111_110011100000001101001001100000
q_pos = 1000
q_neg = 0100

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_101001111010100111010011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_111101000101110011000000000000
w_sum_translation[4] = 000_101001111010100111010011000000
w_carry_translation[4] = 110_111101000101110011000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	111_110011100000001101001001100000 +
	000_000000000000000000000000000000
) = 2 * 111_110011100000001101001001100000 = 
111_100111000000011010010011000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
001_010011110101001110100110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
101_111010001011100110000000000000
w_sum_translation[5] = 111_010011110101001110100110000000
w_carry_translation[5] = 111_111010001011100110000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 11_11 -> q[6] = -1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	111_100111000000011010010011000000 +
	000_000000000000000000000000000000
) = 2 * 111_100111000000011010010011000000 = 
111_001110000000110100100110000000
q_pos = 1000_00
q_neg = 0100_01

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
011_010101110101111001010100000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_001100010100011000010000000000
w_sum_translation[6] = 001_010101110101111001010100000000
w_carry_translation[6] = 111_001100010100011000010000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_11 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	111_001110000000110100100110000000 +
	001_000011000100010100001100000000
) = 2 * 000_010001000101001000110010000000 = 
000_100010001010010001100100000000
q_pos = 1000_000
q_neg = 0100_010

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_101011101011110010101000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
110_011000101000110000100000000000
w_sum_translation[7] = 000_101011101011110010101000000000
w_carry_translation[7] = 000_011000101000110000100000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_00 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_100010001010010001100100000000 +
	000_000000000000000000000000000000
) = 2 * 000_100010001010010001100100000000 = 
001_000100010100100011001000000000
q_pos = 1000_0001
q_neg = 0100_0100

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	001_000100010100100011001000000000 +
	110_111100111011101011110100000000
) = 2 * 000_000001010000001110111100000000 = 
000_000010100000011101111000000000


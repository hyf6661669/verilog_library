参考:
LOW-POWER RADIX-8 DIVIDER, Alberto Nannarelli and Tomas Lang



// ---------------------------------------------------------------------------------------------------------------------------------------
For Radix-8 SRT:
N = log2(8) = 3
进行R8 SRT迭代时, 需要:
1 + WIDTH + 1 + 2 = 32-bit
来表示"w_sum/w_carry", 其中1-bit是符号位, 1-bit是为了做右移操作的位, 2-bit是初始化的时候要将Dividend右移2位的操作
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110100001110011100100011 = 13690659
D[WIDTH-1:0] = 0000000001001001110111011100 = 302556
Q[WIDTH-1:0] = X / D = 45 = 0000000000000000000000101101
REM[WIDTH-1:0] = 13690659 - 302556 * 45 = 75639 = 0000000000010010011101110111

CLZ_X = 4
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 5
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (6 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(7 / 2) = 4;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 1101000011100111001000110000
Divisor[WIDTH-1:0] 		= 1001001110111011100000000000





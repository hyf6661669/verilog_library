// 参考: Radix-64 Floating-Point Divider, Javier D. Bruguera, ARM Austin Design Center

// 为简单起见，仅考虑TABLE I中的第一行，即divisor = 0.1000...., M = 2
// Take FP16 as example..
// for fp16, rem should be 17-bit

a = 0.11010000100
b = 0.10001111111
a / b = 1.01110010111111010001101111001101010010100001000010...
a_scaled = a << 1 = 1.10100001000000
b_scaled = b << 1 = 1.00011111110000

d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000

// ==================================================================================================
rem_init = 00001101000010000
rem_s[0] = rem_init = 00001101000010000
rem_c[0] = 00000000000000000
rem[0] = 00001101000010000

// ================
// BigIter[0]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[0][14:9] + rem_c[0][14:9] = 
001101 + 
000000 = 
001101, belongs to "[13/8, 31/8]" -> q[0] = +2
q_pos = 10
q_neg = 00
q_pos - q_neg = 10

// stage[1]
rem_s[1] = csa(4 * rem_s[0], 4 * rem_c[0], -q[0] * d).s = 10001100001011111
rem_c[1] = csa(4 * rem_s[0], 4 * rem_c[0], -q[0] * d).c = 01100000000000001
-> 
rem[1] = 
00110100001000000 + 
10111000000100000 = 
11101100001100000

rem_s[1][14:9] + rem_c[1][14:9] = 
001100 + 
100000 = 
101100, belongs to "[-32/8, -14/8]" -> q[1] = -2
q_pos = 1000
q_neg = 0010
q_pos - q_neg = 0110

adder_9b = (rem_s[1] << 2)[16:8] + (rem_c[1] << 2)[16:8] = 
001100001 + 
100000000 =
101100001
adder_9b[8:3] = 101100, belongs to "[-32/8, -14/8]" -> q[1] = -2

// stage[2]
rem_s[2] = csa(4 * rem_s[1], 4 * rem_c[1], -q[1] * d).s = 11110111010011000
rem_c[2] = csa(4 * rem_s[1], 4 * rem_c[1], -q[1] * d).c = 00000001011001000
->
rem[2] = 
10110000110000000 + 
01000111111100000 = 
11111000101100000

rem_s[2][14:9] + rem_c[2][14:9] = 
110111 + 
000001 = 
111000, belongs to "[-12/8, -5/8]" -> q[2] = -1
q_pos = 100000
q_neg = 001001
q_pos - q_neg = 010111
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[1] * d) << 2)[16:10] + adder_9b[6:0]
0001111 +
1100001 = 
1110000, adder_7b[6:1] = 111000, belongs to "[-12/8, -4/8]" -> q[2] = -1

// ================
// BigIter[1]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[3] = csa(4 * rem_s[2], 4 * rem_c[2], -q[2] * d).s = 11111011010110000
rem_c[3] = csa(4 * rem_s[2], 4 * rem_c[2], -q[2] * d).c = 00001011011000000
->
rem[3] = 
11100010110000000 + 
00100011111110000 = 
00000110101110000

rem_s[3][14:9] + rem_c[3][14:9] = 
111011 + 
001011 = 
000110, belongs to "[4/8, 12/8]" -> q[3] = +1
q_pos = 10000001
q_neg = 00100100
q_pos - q_neg = 01011101
a / b = 1.0111001011111101000110111100110......

// stage[1]
rem_s[4] = csa(4 * rem_s[3], 4 * rem_c[3], -q[3] * d).s = 00011100111001111
rem_c[4] = csa(4 * rem_s[3], 4 * rem_c[3], -q[3] * d).c = 11011010000000001
->
rem[4] = 
00011010111000000 + 
11011100000010000 = 
11110110111010000

rem_s[4][14:9] + rem_c[4][14:9] = 
011100 + 
011010 = 
110110, belongs to "[-12/8, -5/8]" -> q[4] = -1
q_pos = 1000000100
q_neg = 0010010001
q_pos - q_neg = 0101110011
a / b = 1.0111001011111101000110111100110......

adder_9b = (rem_s[4] << 2)[16:8] + (rem_c[4] << 2)[16:8] = 
011100111 + 
011010000 =
110110111
adder_9b[8:3] = 110110, belongs to "[-12/8, -5/8]" -> q[4] = -1

// stage[2]
rem_s[5] = csa(4 * rem_s[4], 4 * rem_c[4], -q[4] * d).s = 00111000011001000
rem_c[5] = csa(4 * rem_s[4], 4 * rem_c[4], -q[4] * d).c = 11000111001101000
->
rem[5] = 
11011011101000000 + 
00100011111110000 = 
11111111100110000

rem_s[5][14:9] + rem_c[5][14:9] = 
111000 + 
000111 = 
111111, belongs to "[-3/8, 2/8]" -> q[5] = 0
q_pos = 100000010000
q_neg = 001001000100
q_pos - q_neg = 010111001100
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[4] * d) << 2)[16:10] + adder_9b[6:0]
1000111 +
0110111 = 
1111110, adder_7b[6:1] = 111111, belongs to "[-3/8, 3/8]" -> q[5] = 0

// ================
// BigIter[2]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[6] = csa(4 * rem_s[5], 4 * rem_c[5], -q[5] * d).s = 11100001100100000
rem_c[6] = csa(4 * rem_s[5], 4 * rem_c[5], -q[5] * d).c = 00011100110100000
->
rem[6] = 
11111110011000000 + 
00000000000000000 = 
11111110011000000

rem_s[6][14:9] + rem_c[6][14:9] =
100001 + 
011100 = 
111101, belongs to "[-3/8, 3/8]" -> q[6] = 0
q_pos = 10000001000000
q_neg = 00100100010000
q_pos - q_neg = 01011100110000
a / b = 1.0111001011111101000110111100110......

// stage[1]
rem_s[7] = csa(4 * rem_s[6], 4 * rem_c[6], -q[6] * d).s = 10000110010000000
rem_c[7] = csa(4 * rem_s[6], 4 * rem_c[6], -q[6] * d).c = 01110011010000000
->
rem[7] = 
11111001100000000 + 
00000000000000000 = 
11111001100000000

rem_s[7][14:9] + rem_c[7][14:9] = 
000110 + 
110011 = 
111001, belongs to "[-12/8, -4/8]" -> q[7] = -1
q_pos = 1000000100000000
q_neg = 0010010001000001
q_pos - q_neg = 0101110010111111
a / b = 1.0111001011111101000110111100110......

adder_9b = (rem_s[7] << 2)[16:8] + (rem_c[7] << 2)[16:8] = 
000110010 + 
110011010 =
111001100
adder_9b[8:3] = 111001, belongs to "[-12/8, -5/8]" -> q[7] = -1

// stage[2]
rem_s[8] = csa(4 * rem_s[7], 4 * rem_c[7], -q[7] * d).s = 11110111111110000
rem_c[8] = csa(4 * rem_s[7], 4 * rem_c[7], -q[7] * d).c = 00010010000000000
->
rem[8] = 
11100110000000000 + 
00100011111110000 = 
00001001111110000

rem_s[8][14:9] + rem_c[8][14:9] = 
110111 + 
010010 = 
001001, belongs to "[4/8, 11/8]" -> q[8] = +1
q_pos = 100000010000000001
q_neg = 001001000100000100
q_pos - q_neg = 010111001011111101
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[7] * d) << 2)[16:10] + adder_9b[6:0]
1000111 +
1001100 = 
0010011, adder_7b[6:1] = 001001, belongs to "[4/8, 12/8]" -> q[8] = +1

// ================
// BigIter[3]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[9] = csa(4 * rem_s[8], 4 * rem_c[8], -q[8] * d).s = 01001011111001111
rem_c[9] = csa(4 * rem_s[8], 4 * rem_c[8], -q[8] * d).c = 10111000000000001
->
rem[9] = 
00100111111000000 + 
11011100000010000 = 
00000011111010000

rem_s[9][14:9] + rem_c[9][14:9] =
001011 + 
111000 = 
000011, belongs to "[-3/8, 3/8]" -> q[9] = 0
q_pos = 10000001000000000100
q_neg = 00100100010000010000
q_pos - q_neg = 01011100101111110100
a / b = 1.0111001011111101000110111100110......

// stage[1]
rem_s[10] = csa(4 * rem_s[9], 4 * rem_c[9], -q[9] * d).s = 00101111100111100
rem_c[10] = csa(4 * rem_s[9], 4 * rem_c[9], -q[9] * d).c = 11100000000000100
->
rem[10] = 
00001111101000000 + 
00000000000000000 = 
00001111101000000

rem_s[10][14:9] + rem_c[10][14:9] = 
101111 + 
100000 = 
001111, belongs to "[13/8, 31/8]" -> q[10] = +2
q_pos = 1000000100000000010010
q_neg = 0010010001000001000000
q_pos - q_neg = 0101110010111111010010
a / b = 1.0111001011111101000110111100110......

adder_9b = (rem_s[10] << 2)[16:8] + (rem_c[10] << 2)[16:8] = 
101111100 + 
100000000 =
001111100
adder_9b[8:3] = 001111, belongs to "[13/8, 30/8]" -> q[10] = +2

// stage[2]
rem_s[11] = csa(4 * rem_s[10], 4 * rem_c[10], -q[10] * d).s = 10000110011111111
rem_c[11] = csa(4 * rem_s[10], 4 * rem_c[10], -q[10] * d).c = 01110000000100001
->
rem[11] = 
00111110100000000 + 
10111000000100000 = 
11110110100100000

rem_s[11][14:9] + rem_c[11][14:9] = 
000110 + 
110000 = 
110110, belongs to "[-12/8, -4/8]" -> q[11] = -1
q_pos = 100000010000000001001000
q_neg = 001001000100000100000001
q_pos - q_neg = 010111001011111101000111
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[10] * d) << 2)[16:10] + adder_9b[6:0]
1110000 +
1111100 = 
1101100, adder_7b[6:1] = 110110, belongs to "[-12/8, -5/8]" -> q[11] = -1

// ================
// BigIter[4]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[12] = 11111010010001000
rem_c[12] = 00000011111101000
->
rem[12] = 
11011010010000000 + 
00100011111110000 = 
11111110001110000

rem_s[12][14:9] + rem_c[12][14:9] =
111010 + 
000011 = 
111101, belongs to "[-3/8, 3/8]" -> q[12] = 0
q_pos = 10000001000000000100100000
q_neg = 00100100010000010000000100
q_pos - q_neg = 01011100101111110100011100
a / b = 1.0111001011111101000110111100110......

// stage[1]
rem_s[13] = 11101001000100000
rem_c[13] = 00001111110100000
->
rem[13] = 
11111000111000000 + 
00000000000000000 = 
11111000111000000

rem_s[13][14:9] + rem_c[13][14:9] = 
101001 + 
001111 = 
111000, belongs to "[-12/8, -4/8]" -> q[13] = -1
q_pos = 1000000100000000010010000000
q_neg = 0010010001000001000000010001
q_pos - q_neg = 0101110010111111010001101111
1.01110010111111010001101111001101010010100001000010...

adder_9b = (rem_s[13] << 2)[16:8] + (rem_c[13] << 2)[16:8] = 
101001000 + 
001111110 =
111000110
adder_9b[8:3] = 111000, belongs to "[-12/8, -5/8]" -> q[13] = -1

// stage[2]
rem_s[14] = 10111000111110000
rem_c[14] = 01001110100000000
->
rem[14] = 
11100011100000000 + 
00100011111110000 = 
00000111011110000

rem_s[14][14:9] + rem_c[14][14:9] = 
111000 + 
001110 = 
000110, belongs to "[4/8, 12/8]" -> q[14] = +1
q_pos = 100000010000000001001000000001
q_neg = 001001000100000100000001000100
q_pos - q_neg = 010111001011111101000110111101
1.01110010111111010001101111001101010010100001000010...

adder_7b = ((-q[13] * d) << 2)[16:10] + adder_9b[6:0]
1000111 +
1000110 = 
0001101, adder_7b[6:1] = 000110, belongs to "[4/8, 12/8]" -> q[14] = +1

// ================
// BigIter[5]
d   = 00100011111110000
2d  = 01000111111100000
~d  = 11011100000001111
~2d = 10111000000011111
-d  = 11011100000010000
-2d = 10111000000100000
// ================
// stage[0]
rem_s[15] = 00000101111001111
rem_c[15] = 11110100000000001
->
rem[15] = 
00011101111000000 + 
11011100000010000 = 
11111001111010000

rem_s[15][14:9] + rem_c[15][14:9] =
000101 + 
110100 = 
111001, belongs to "[-12/8, -4/8]" -> q[15] = -1
q_pos = 10000001000000000100100000000100
q_neg = 00100100010000010000000100010001
q_pos - q_neg = 01011100101111110100011011110011
1.01110010111111010001101111001101010010100001000010...

// TODO
// stage[1]
rem_s[13] = 11101001000100000
rem_c[13] = 00001111110100000
->
rem[13] = 
11111000111000000 + 
00000000000000000 = 
11111000111000000

rem_s[13][14:9] + rem_c[13][14:9] = 
101001 + 
001111 = 
111000, belongs to "[-12/8, -4/8]" -> q[13] = -1
q_pos = 1000000100000000010010000000
q_neg = 0010010001000001000000010001
q_pos - q_neg = 0101110010111111010001101111
1.01110010111111010001101111001101010010100001000010...

adder_9b = (rem_s[13] << 2)[16:8] + (rem_c[13] << 2)[16:8] = 
101001000 + 
001111110 =
111000110
adder_9b[8:3] = 111000, belongs to "[-12/8, -5/8]" -> q[13] = -1

// stage[2]
rem_s[14] = 10111000111110000
rem_c[14] = 01001110100000000
->
rem[14] = 
11100011100000000 + 
00100011111110000 = 
00000111011110000

rem_s[14][14:9] + rem_c[14][14:9] = 
111000 + 
001110 = 
000110, belongs to "[4/8, 12/8]" -> q[14] = +1
q_pos = 100000010000000001001000000001
q_neg = 001001000100000100000001000100
q_pos - q_neg = 010111001011111101000110111101
1.01110010111111010001101111001101010010100001000010...

adder_7b = ((-q[13] * d) << 2)[16:10] + adder_9b[6:0]
1000111 +
1000110 = 
0001101, adder_7b[6:1] = 000110, belongs to "[4/8, 12/8]" -> q[14] = +1







测试Radix-2 fpsqrt

// ---------------------------------------------------------------------------------------------------------------------------------------
fp16
// ---------------------------------------------------------------------------------------------------------------------------------------
X[11-1:0] = 1.1010_0011_00 = 1.636718750
X[11] = 0
sqrt(X[11:0]) = 1.27934309315367001749873265846519061894120987869294 = 1.0100011110_0_0001...


stage[0]:
X[11:10] - 01 = 
01 - 
01 = 
{0_00} >= 0
rem[0] = 00
q[11] = 1

stage[1]:
{rem[0][1:0], X[9:8]} - {0, q[11], 01}
0010 -
0101 = 
{1_1101} < 0
rem[1] = 010
q[11:10] = 10

stage[2]:
{rem[1][2:0], X[7:6]} - {0, q[11:10], 01}
01010 -
01001 = 
{0_00001} >= 0
rem[2] = 0001
q[11:9] = 101

stage[3]:
{rem[2][3:0], X[5:4]} - {0, q[11:9], 01}
000100 -
010101 = 
{1_101111} < 0
rem[3] = 00100
q[11:8] = 1010

stage[4]:
{rem[3][4:0], X[3:2]} - {0, q[11:8], 01}
0010011 -
0101001 = 
{1_1101010} < 0
rem[4] = 010011
q[11:7] = 10100

stage[5]:
{rem[4][5:0], X[1:0]} - {0, q[11:7], 01}
01001100 -
01010001 = 
{1_11111011} < 0
rem[5] = 1001100
q[11:6] = 101000

stage[6]:
{rem[5][6:0], 00} - {0, q[11:6], 01}
100110000 -
010100001 = 
{0_010001111} >= 0
rem[6] = 10001111
q[11:5] = 1010001

stage[7]:
{rem[6][7:0], 00} - {0, q[11:5], 01}
1000111100 -
0101000101 = 
{0_0011110111} >= 0
rem[7] = 011110111
q[11:4] = 10100011

stage[8]:
{rem[7][8:0], 00} - {0, q[11:4], 01}
01111011100 -
01010001101 = 
{0_00101001111} >= 0
rem[8] = 0101001111
q[11:3] = 101000111

stage[9]:
{rem[8][9:0], 00} - {0, q[11:3], 01}
010100111100 -
010100011101 = 
{0_000000011111} >= 0
rem[9] = 00000011111
q[11:2] = 1010001111

stage[10]:
{rem[9][10:0], 00} - {0, q[11:2], 01}
0000001111100 -
0101000111101 = 
{1_1011000111111} < 0
rem[10] = 000001111100
q[11:1] = 10100011110

stage[11]:
{rem[10][11:0], 00} - {0, q[11:1], 01}
00000111110000 -
01010001111001 = 
{1_10110101110111} < 0
rem[11] = 0000111110000
q[11:0] = 101000111100


// ---------------------------------------------------------------------------------------------------------------------------------------
X[11-1:0] = 1.1010_0011_00
X[12-1:0] << 1 = 11.0100_0110_00 = 3.27343750
sqrt(X[12-1:0]) = 1.1100111100_1_0101111110...

1.11001111001 ^ 2 = 11.0100010111010100110001
11.0100011000 - 11.0100010111010100110001 = 0.0000000000101011001111


stage[0]:
X[11:10] - 01 = 
11 - 
01 = 
{0_10} >= 0
rem[0] = 10
q[11] = 1

stage[1]:
{rem[0][1:0], X[9:8]} - {0, q[11], 01}
1001 -
0101 = 
{0_100} >= 0
rem[1] = 100
q[11:10] = 11

stage[2]:
{rem[1][2:0], X[7:6]} - {0, q[11:10], 01}
10000 -
01101 = 
{0_00011} >= 0
rem[2] = 0011
q[11:9] = 111

stage[3]:
{rem[2][3:0], X[5:4]} - {0, q[11:9], 01}
001101 -
011101 = 
{1_110000} < 0
rem[3] = 01101
q[11:8] = 1110

stage[4]:
{rem[3][4:0], X[3:2]} - {0, q[11:8], 01}
0110110 -
0111001 = 
{1_1111101} < 0
rem[4] = 110110
q[11:7] = 11100

stage[5]:
{rem[4][5:0], X[1:0]} - {0, q[11:7], 01}
11011000 -
01110001 = 
{0_01100111} >= 0
rem[5] = 1100111
q[11:6] = 111001

stage[6]:
{rem[5][6:0], 00} - {0, q[11:6], 01}
110011100 -
011100101 = 
{0_010110111} >= 0
rem[6] = 10110111
q[11:5] = 1110011

stage[7]:
{rem[6][7:0], 00} - {0, q[11:5], 01}
1011011100 -
0111001101 = 
{0_0100001111} >= 0
rem[7] = 100001111
q[11:4] = 11100111

stage[8]:
{rem[7][8:0], 00} - {0, q[11:4], 01}
10000111100 -
01110011101 = 
{0_00010011111} >= 0
rem[8] = 0010011111
q[11:3] = 111001111

stage[9]:
{rem[8][9:0], 00} - {0, q[11:3], 01}
001001111100 -
011100111101 = 
{1_101100111111} < 0
rem[9] = 01001111100
q[11:2] = 1110011110

stage[10]:
{rem[9][10:0], 00} - {0, q[11:2], 01}
0100111110000 -
0111001111001 = 
{1_1101101110111} < 0
rem[10] = 100111110000
q[11:1] = 11100111100

stage[11]:
{rem[10][11:0], 00} - {0, q[11:1], 01}
10011111000000 -
01110011110001 = 
{0_00101011001111} >= 0
rem[11] = 0101011001111
q[11:0] = 111001111001

// ========================================================================
由上述计算实例可知，为得到"N-bit"的root, 需要使用"(N + 2)-bit"的全加器，再将符号位考虑进来，则需要"(N + 3)-bit"的全加器



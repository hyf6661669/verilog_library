保持divisor不动，将dividend右移"CLZ_DIFF = CLZ_D - CLZ_X"使得2者的MSB对齐，注意需要使用寄存器记录dividend右移出去的那些数字
然后按照SRT的结果来迭代计算每一步的余数，在迭代结束的时候这个数据通路得到的REM结果就直接是最终的REM结果，不需要额外的右移操作.
相当于把后处理中的右移放在前处理完成了

设:
WIDTH = 28
REM_W = 1 + (2 * WIDTH) + 3 = 60

X[WIDTH-1:0] = 1000010110011111011100111011 = 140113723
D[WIDTH-1:0] = 0000000000000110000001000011 = 24643
Q[WIDTH-1:0] = X / D = 5685 = 0000000000000001011000110101
REM[WIDTH-1:0] = 140113723 - 24643 * 5685 = 18268 = 0000000000000100011101011100

CLZ_X = 0
CLZ_D = 13
CLZ_DIFF = CLZ_D - CLZ_X = 13
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (14 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(15 / 2) = 8;

+ D = 0_00000000000001100000010000110000000000000000000000000000000
+2D = 0_00000000000011000000100001100000000000000000000000000000000
- D = 1_11111111111110011111101111010000000000000000000000000000000
-2D = 1_11111111111100111111011110100000000000000000000000000000000


X >> (CLZ_DIFF + 2 + r_shift_num) = 0_00000000000000001000010110011111011100111011000000000000000
w[0] = 0_00000000000000001000010110011111011100111011000000000000000

q[1] = 0
w[1] = 4 * w[0] - q[1] * D = 
0_00000000000000100001011001111101110011101100000000000000000 + 
0_00000000000000000000000000000000000000000000000000000000000 = 
0_00000000000000100001011001111101110011101100000000000000000

q[2] = +1
w[2] = 4 * w[1] - q[2] * D = 
0_00000000000010000101100111110111001110110000000000000000000 + 
1_11111111111110011111101111010000000000000000000000000000000 = 
0_00000000000000100101010111000111001110110000000000000000000

q[3] = +2
w[3] = 4 * w[2] - q[3] * D = 
0_00000000000010010101011100011100111011000000000000000000000 + 
1_11111111111100111111011110100000000000000000000000000000000 = 
1_11111111111111010100111010111100111011000000000000000000000

q[4] = -2
w[4] = 4 * w[3] - q[4] * D = 
1_11111111111101010011101011110011101100000000000000000000000 + 
0_00000000000011000000100001100000000000000000000000000000000 = 
0_00000000000000010100001101010011101100000000000000000000000

q[5] = +1
w[5] = 4 * w[4] - q[5] * D = 
0_00000000000001010000110101001110110000000000000000000000000 + 
1_11111111111110011111101111010000000000000000000000000000000 = 
1_11111111111111110000100100011110110000000000000000000000000

q[6] = -1
w[6] = 4 * w[5] - q[6] * D = 
1_11111111111111000010010001111011000000000000000000000000000 + 
0_00000000000001100000010000110000000000000000000000000000000 = 
0_00000000000000100010100010101011000000000000000000000000000

q[7] = +1
w[7] = 4 * w[6] - q[7] * D = 
0_00000000000010001010001010101100000000000000000000000000000 + 
1_11111111111110011111101111010000000000000000000000000000000 = 
0_00000000000000101001111001111100000000000000000000000000000

q[8] = +2
w[8] = 4 * w[7] - q[8] * D = 
0_00000000000010100111100111110000000000000000000000000000000 + 
1_11111111111100111111011110100000000000000000000000000000000 = 
1_11111111111111100111000110010000000000000000000000000000000

w[8] + D = 
1_11111111111111100111000110010000000000000000000000000000000 + 
0_00000000000001100000010000110000000000000000000000000000000 = 
0_00000000000001000111010111000000000000000000000000000000000









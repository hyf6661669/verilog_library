接"test_broken_1.sv".
在之前的通过overlap多个Radix-2以得到"High-Radix的"例子中，发现如果迭代开始时没有把"Dividend"规格化到区间"[1, 2)", 
会遇到很多原来不会出现的问题。
初步分析是因为前处理操作中如果没有将"Dividend"规格化到区间"[1, 2)", 则前面的几个bit的商应当是0, 但是按照paper给出的商选择函数来计算, 会选择出非0的商, 
这导致最后的结果出错。


那么尝试在前处理步骤中不再将"Dividend"右移了, 而是在最后一次大迭代计算中改变商的选择函数以及余数的计算方式，
从而生成正确的商和余数。
这样也不用增加迭代过程中"w_sum[i]/w_carry[i]"的宽度了.
// ---------------------------------------------------------------------------------------------------------------------------------------
Radix-8:
iter_num % 3 =
0: 最后一次大迭代的第2次小迭代计算出的结果刚好是最终的商，无需改变"1 ~ 2"次的小迭代中的商选择函数和余数的计算方式;
1: 最后一次大迭代的第0次小迭代计算出的结果刚好是最终的商，需要改变"1 ~ 2"次的小迭代中的商选择函数和余数的计算方式, 强制:
q_modified[2] = q_modified[1] = 0;
w_sum_modified[2] = w_sum_modified[1] = w_sum[0];
w_carry_modified[2] = w_carry_modified[1] = w_carry[0];
2: 最后一次大迭代的第1次小迭代计算出的结果刚好是最终的商，需要改变"2"次的小迭代中的商选择函数和余数的计算方式, 强制:
q_modified[2] = 0;
w_sum_modified[2] = w_sum[1];
w_carry_modified[2] = w_carry[1];
// ---------------------------------------------------------------------------------------------------------------------------------------
Radix-16:
iter_num % 4 =
0: 最后一次大迭代的第3次小迭代计算出的结果刚好是最终的商，无需改变"1 ~ 3"次的小迭代中的商选择函数和余数的计算方式;
1: 最后一次大迭代的第0次小迭代计算出的结果刚好是最终的商，需要改变"1 ~ 3"次的小迭代中的商选择函数和余数的计算方式, 强制:
q_modified[3] = q_modified[2] = q_modified[1] = 0;
w_sum_modified[3] = w_sum_modified[2] = w_sum_modified[1] = w_sum[0];
w_carry_modified[3] = w_carry_modified[2] = w_carry_modified[1] = w_carry[0];
2: 最后一次大迭代的第1次小迭代计算出的结果刚好是最终的商，需要改变"2 ~ 3"次的小迭代中的商选择函数和余数的计算方式, 强制:
q_modified[3] = q_modified[2] = 0;
w_sum_modified[3] = w_sum_modified[2] = w_sum[1];
w_carry_modified[3] = w_carry_modified[2] = w_carry[1];
3: 最后一次大迭代的第2次小迭代计算出的结果刚好是最终的商，需要改变"3"次的小迭代中的商选择函数和余数的计算方式, 强制:
q_modified[3] = 0;
w_sum_modified[3] = w_sum[2];
w_carry_modified[3] = w_carry[2];

这样又有新的问题，即现在一次大迭代中的所有小迭代都可能是最后一次迭代，而我们又为最后一次迭代使用了特殊的QDS(详见"division_test6.sv").
那么对于每次大迭代中的第"0"次小迭代来说, QDS会变慢一点，因为其要受到上次大迭代中最后一次小迭代的商数字的影响(寄存器输出), 对于第"1 ~ (N-1)"次小迭代来说, QDS并不会变慢，
因为它们的QDS由上一次小迭代的商数字以及"iter_num_last"决定，而上一次小迭代的商数字计算出来之后，还要经过"Mux"操作才能得到下一次小迭代的"w_sum[i]/w_carry[i]".
那么在"Mux"的同时也可以确定出下一次小迭代的QDS.

或者可以仿照ARM的作法, 在每次大迭代的末尾根据"iter_num_last"的值进行"MUX"操作, 似乎各有优劣...



// ---------------------------------------------------------------------------------------------------------------------------------------
在后处理的时候，将"q_pos/q_neg"右移几位之后再计算"q_calculated", 设"iter_num_last"为最后一次大迭代步骤中记录还需要几次小迭代的计数器.
// ---------------------------------------------------------------------------------------------------------------------------------------
Radix-8:
iter_num_last = 1, 2, 3;
r_shift_num = 3 - iter_num_last -> 
iter_num_last = 1, r_shift_num = 2;
iter_num_last = 2, r_shift_num = 1;
iter_num_last = 3, r_shift_num = 0;
// ---------------------------------------------------------------------------------------------------------------------------------------
Radix-16:
iter_num_last = 1, 2, 3, 4;
r_shift_num = 4 - iter_num_last -> 
iter_num_last = 1, r_shift_num = 3;
iter_num_last = 2, r_shift_num = 2;
iter_num_last = 3, r_shift_num = 1;
iter_num_last = 4, r_shift_num = 0;
// ---------------------------------------------------------------------------------------------------------------------------------------
下面搞几个测试来看看.
WIDTH = 28;
将3个Radix-2串联起来形成Radix-8算法, 即:
N = 8;
(WIDTH + 1 + log2(N)) = 32;

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000000010100010100001100001 = 665697
D[WIDTH-1:0] = 0000000000010011100001111111 = 79999
Q[WIDTH-1:0] = X / D = 8 = 0000000000000000000000001000
REM[WIDTH-1:0] = 1189985 - 79999 * 8 = 25705 = 0000000000000110010001101001

CLZ_X = 8
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 3
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(5 / 3) = 2;
iter_num_last = 2;
r_shift_num = 3 - iter_num_last = 1;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1010001010000110000100000000
Divisor[WIDTH-1:0] 		= 1001110000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_001110000111111100000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_011100001111111000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_110001111000000100000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_100011110000001000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[3 * iter_num - r_shift_num] = w[5] = 111_001000001010011000000000000 < 0
// 最后一次迭代的商
q[final] = q[3 * iter_num - r_shift_num] = q[5] = -1;
q_pos = 1001_00 >> r_shift_num = 10010
q_neg = 0000_10 >> r_shift_num = 00001
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 00010001
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0001000
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 2)[0 +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1100100000101001100000000000 + 1001110000111111100000000000 = 
0110010001101001000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0110010001101001000000000000 >> 11 = 
0000000000000110010001101001

q[4] = +1
q[5] = -1
w[5] = 111_001000001010011000000000000 < 0
w[5] / 2 = 111_100100000101001100000000000
111_100100000101001100000000000 + D = 
111_100100000101001100000000000 + 001_001110000111111100000000000 = 
000_110010001101001000000000000

0110010001101001000000000000 >> (CLZ_D + 1) = 
0000000000000110010001101001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_010001010000110000100000000
w_sum_translation[0] = w_sum[0] =  001_010001010000110000100000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 2){1'b0}} = 000_000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_100010100001100001000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_100011110000001000000000000
w_sum_translation[1] = 000_100010100001100001000000000
w_carry_translation[1] = 111_100011110000001000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_010001010000110000100000000 +
	110_110001111000000100000000000
) = 2 * 000_000011001000110100100000000 = 
000_000110010001101001000000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_000101000011000010000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_000111100000010000000000000
w_sum_translation[2] = 001_000101000011000010000000000
w_carry_translation[2] = 111_000111100000010000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_000110010001101001000000000 +
	000_000000000000000000000000000
) = 2 * 000_000110010001101001000000000 = 
000_001100100011010010000000000
q_pos = 100
q_neg = 000

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_001010000110000100000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_001111000000100000000000000
w_sum_translation[3] = 000_001010000110000100000000000
w_carry_translation[3] = 000_001111000000100000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_00 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_001100100011010010000000000 +
	000_000000000000000000000000000
) = 2 * 000_001100100011010010000000000 = 
000_011001000110100100000000000
q_pos = 1001
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
101_101001111101000000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_101100000000010000000000000
w_sum_translation[4] = 111_101001111101000000000000000
w_carry_translation[4] = 110_101100000000010000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_10 -> q[5] = -1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_011001000110100100000000000 +
	110_110001111000000100000000000
) = 2 * 111_001010111110101000000000000 = 
110_010101111101010000000000000
q_pos = 1001_0
q_neg = 0000_1

// 需要修改这个小迭代开始后面的的商和余数的生成逻辑
q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	110_010101111101010000000000000 +
	001_001110000111111100000000000
) = 2 * 111_100100000101001100000000000 = 
111_001000001010011000000000000
q_pos = 1001_00
q_neg = 0000_10
w[6] = w[5] = 111_001000001010011000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000001000001011111100000010 = 2146050
D[WIDTH-1:0] = 0000000000010000100001111111 = 67711
Q[WIDTH-1:0] = X / D = 31 = 0000000000000000000000011111
REM[WIDTH-1:0] = 2146050 - 67711 * 31 = 47009 = 0000000000001011011110100001

CLZ_X = 6
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 5
迭代次数
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(7 / 3) = 3;
iter_num_last = 1;
r_shift_num = 3 - iter_num_last = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000001011111100000010000000
Divisor[WIDTH-1:0] 		= 1000010000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_000010000111111100000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_000100001111111000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_111101111000000100000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_111011110000001000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// TODO
// 最后一次迭代的余数
w[final] = w[3 * iter_num - r_shift_num] = w[7] = 000_110011011000011000000000000 >= 0
// 最后一次迭代的商
q[final] = q[3 * iter_num - r_shift_num] = q[7] = -1;
q_pos = 1000_000
q_neg = 0000_001
q_calculated_pre[(WIDTH + 1) - 1:0] = q_pos[(WIDTH + 1) - 1:0] - q_neg[(WIDTH + 1) - 1:0] = 00111111
q_calculated[WIDTH-1:0] = (q_calculated_pre[(WIDTH + 1) - 1:0] - (w[final] < 0))[WIDTH:1] = 0011111
remainder_calculated_pre[WIDTH-1:0] = ((w[final] / 4)[log2(N) +: WIDTH] + (w[final] < 0 ? Divisor : {(WIDTH){1'b0}}))[WIDTH-1:0] = 
1101011110010001000000000000 + 1000010000111111100000000000 = 
0101101111010000100000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
0101101111010000100000000000 >> 11 = 
0000000000001011011110100001
// 结果正确
// TEST
w[7] / 2 = 0011001101100001100000000000
0011001101100001100000000000 + (D) = 
0011001101100001100000000000 + 1000010000111111100000000000 = 
1011011110100001000000000000

1011011110100001000000000000 >> (CLZ_D + 1) = 
0000000000001011011110100001

// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_000001011111100000010000000
w_sum_translation[0] = w_sum[0] =  001_000001011111100000010000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
010_000010111111000000100000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_111011110000001000000000000
w_sum_translation[1] = 000_000010111111000000100000000
w_carry_translation[1] = 111_111011110000001000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 00_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_000001011111100000010000000 +
	110_111101111000000100000000000
) = 2 * 111_111111010111100100010000000 = 
111_111110101111001000100000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_000101111110000001000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_110111100000010000000000000
w_sum_translation[2] = 000_000101111110000001000000000
w_carry_translation[2] = 111_110111100000010000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	111_111110101111001000100000000 +
	000_000000000000000000000000000
) = 2 * 111_111110101111001000100000000 = 
111_111101011110010001000000000
q_pos = 100
q_neg = 000

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_001011111100000010000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_101111000000100000000000000
w_sum_translation[3] = 000_001011111100000010000000000
w_carry_translation[3] = 111_101111000000100000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	111_111101011110010001000000000 +
	000_000000000000000000000000000
) = 2 * 111_111101011110010001000000000 = 
111_111010111100100010000000000
q_pos = 1000
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_010111111000000100000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_011110000001000000000000000
w_sum_translation[4] = 000_010111111000000100000000000
w_carry_translation[4] = 111_011110000001000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_11 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	111_111010111100100010000000000 +
	000_000000000000000000000000000
) = 2 * 111_111010111100100010000000000 = 
111_110101111001000100000000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_101111110000001000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_111100000010000000000000000
w_sum_translation[5] = 000_101111110000001000000000000
w_carry_translation[5] = 110_111100000010000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_10 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	111_110101111001000100000000000 +
	000_000000000000000000000000000
) = 2 * 111_110101111001000100000000000 = 
111_101011110010001000000000000
q_pos = 1000_00
q_neg = 0000_00

// 第3次大迭代
w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_011111100000010000000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_111000000100000000000000000
w_sum_translation[6] = 111_011111100000010000000000000
w_carry_translation[6] = 111_111000000100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 11_11 -> q[7] = -1
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	111_101011110010001000000000000 +
	000_000000000000000000000000000
) = 2 * 111_101011110010001000000000000 = 
111_010111100100010000000000000
q_pos = 1000_000
q_neg = 0000_001

w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	111_010111100100010000000000000 +
	001_000010000111111100000000000
) = 2 * 000_011001101100001100000000000 = 
000_110011011000011000000000000

// 需要修改这个小迭代开始后面的的商和余数的生成逻辑
q[8] = 0
w[8] = w[7];

q[9] = 0
w[9] = w[8];



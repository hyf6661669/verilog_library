测试DW中使用的radix-4 restoring算法, 有符号除法, 求被除数的绝对值.

// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 32;
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 11111010000110010100011010111011 = -99006789
D[WIDTH-1:0] = 11111111111111111111101110111111 = -1089
Q[WIDTH-1:0] = X / D = 90915 = 00000000000000010110001100100011
R[WIDTH-1:0] = -(99006789 - 1089 * 90915) = -354 = 11111111111111111111111010011110
abs(X) = 00000101111001101011100101000101



已知"D < 0"
下面的"X"都是"abs(X)"

radix-2有符号除法的计算过程:
stage[0]:
force_q_to_zero[0] = ~&(D[31:1]) | ~|(D[0:0]) = 1 -> rem[0] = X[31] = 0
q = 0

stage[1]:
force_q_to_zero[1] = ~&(D[31:2]) | ~|(D[1:0]) = 1
{cout[1], sum[1]} = {rem[0], X[30]} + D[1:0] = 
00 + 
11 = 
{0_11} < 0
rem[1] = 00
q = 00

stage[2]:
force_q_to_zero[2] = ~&(D[31:3]) | ~|(D[2:0]) = 1
{cout[2], sum[2]} = {rem[1], X[29]} + D[2:0] = 
000 + 
111 = 
{0_111} < 0
rem[2] = 000
q = 000

stage[3]:
force_q_to_zero[3] = ~&(D[31:4]) | ~|(D[3:0]) = 1
{cout[3], sum[3]} = {rem[2], X[28]} + D[3:0] = 
0000 + 
1111 = 
{0_1111} < 0
rem[3] = 0000
q = 0000

stage[4]:
force_q_to_zero[4] = ~&(D[31:5]) | ~|(D[4:0]) = 1
{cout[4], sum[4]} = {rem[3], X[27]} + D[4:0] = 
00000 + 
11111 = 
{0_11111} < 0
rem[4] = 00000
q = 00000

stage[5]:
force_q_to_zero[5] = ~&(D[31:6]) | ~|(D[5:0]) = 1
{cout[5], sum[5]} = {rem[4], X[26]} + D[5:0] = 
000001 + 
111111 = 
{1_000000} >= 0
rem[5] = 000001
q = 000000

stage[6]:
force_q_to_zero[6] = ~&(D[31:7]) | ~|(D[6:0]) = 1
{cout[6], sum[6]} = {rem[5], X[25]} + D[6:0] = 
0000010 + 
0111111 = 
{0_1000001} < 0
rem[6] = 0000010
q = 0000000

stage[7]:
force_q_to_zero[7] = ~&(D[31:8]) | ~|(D[7:0]) = 1
{cout[7], sum[7]} = {rem[6], X[24]} + D[7:0] = 
00000101 + 
10111111 = 
{0_11000100} < 0
rem[7] = 00000101
q = 00000000

stage[8]:
force_q_to_zero[8] = ~&(D[31:9]) | ~|(D[8:0]) = 1
{cout[8], sum[8]} = {rem[7], X[23]} + D[8:0] = 
000001011 + 
110111111 = 
{0_111001010} < 0
rem[8] = 000001011
q = 000000000

stage[9]:
force_q_to_zero[9] = ~&(D[31:10]) | ~|(D[9:0]) = 1
{cout[9], sum[9]} = {rem[8], X[22]} + D[9:0] = 
0000010111 + 
1110111111 = 
{0_1111010110} < 0
rem[9] = 0000010111
q = 0000000000

stage[10]:
force_q_to_zero[10] = ~&(D[31:11]) | ~|(D[10:0]) = 0
{cout[10], sum[10]} = {rem[9], X[21]} + D[10:0] = 
00000101111 + 
01110111111 = 
{0_01111101110} < 0
rem[10] = 00000101111
q = 00000000000

stage[11]:
force_q_to_zero[11] = ~&(D[31:12]) | ~|(D[11:0]) = 0
{cout[11], sum[11]} = {rem[10], X[20]} + D[11:0] = 
000001011110 + 
101110111111 = 
{0_110000011101} < 0
rem[11] = 000001011110
q = 000000000000

stage[12]:
force_q_to_zero[12] = ~&(D[31:13]) | ~|(D[12:0]) = 0
{cout[12], sum[12]} = {rem[11], X[19]} + D[12:0] = 
0000010111100 + 
1101110111111 = 
{0_1110001111011} < 0
rem[12] = 0000010111100
q = 0000000000000

stage[13]:
force_q_to_zero[13] = ~&(D[31:14]) | ~|(D[13:0]) = 0
{cout[13], sum[13]} = {rem[12], X[18]} + D[13:0] = 
00000101111001 + 
11101110111111 = 
{0_11110100111000} < 0
rem[13] = 00000101111001
q = 00000000000000

stage[14]:
force_q_to_zero[14] = ~&(D[31:15]) | ~|(D[14:0]) = 0
{cout[14], sum[14]} = {rem[13], X[17]} + D[14:0] = 
000001011110011 + 
111101110111111 = 
{0_111111010110010} < 0
rem[14] = 000001011110011
q = 000000000000000

stage[15]:
force_q_to_zero[15] = ~&(D[31:16]) | ~|(D[15:0]) = 0
{cout[15], sum[15]} = {rem[14], X[16]} + D[15:0] = 
0000010111100110 + 
1111101110111111 = 
{1_0000000110100101} >= 0
rem[15] = 0000000110100101
q = 0000000000000001

stage[16]:
force_q_to_zero[16] = ~&(D[31:17]) | ~|(D[16:0]) = 0
{cout[16], sum[16]} = {rem[15], X[15]} + D[16:0] = 
00000001101001011 + 
11111101110111111 = 
{0_11111111100001010} < 0
rem[16] = 00000001101001011
q = 00000000000000010

stage[17]:
force_q_to_zero[17] = ~&(D[31:18]) | ~|(D[17:0]) = 0
{cout[17], sum[17]} = {rem[16], X[14]} + D[17:0] = 
000000011010010110 + 
111111101110111111 = 
{1_000000001001010101} >= 0
rem[17] = 000000001001010101
q = 000000000000000101

stage[18]:
force_q_to_zero[18] = ~&(D[31:19]) | ~|(D[18:0]) = 0
{cout[18], sum[18]} = {rem[17], X[13]} + D[18:0] = 
0000000010010101011 + 
1111111101110111111 = 
{1_0000000000001101010} >= 0
rem[18] = 0000000000001101010
q = 0000000000000001011

stage[19]:
force_q_to_zero[19] = ~&(D[31:20]) | ~|(D[19:0]) = 0
{cout[19], sum[19]} = {rem[18], X[12]} + D[19:0] = 
00000000000011010101 + 
11111111101110111111 = 
{0_11111111110010010100} < 0
rem[19] = 0_00000000000011010101
q = 00000000000000010110

stage[20]:
force_q_to_zero[20] = ~&(D[31:21]) | ~|(D[20:0]) = 0
{cout[20], sum[20]} = {rem[19], X[11]} + D[20:0] = 
000000000000110101011 + 
111111111101110111111 = 
{0_111111111110101101010} < 0
rem[20] = 000000000000110101011
q = 000000000000000101100

stage[21]:
force_q_to_zero[21] = ~&(D[31:22]) | ~|(D[21:0]) = 0
{cout[21], sum[21]} = {rem[20], X[10]} + D[21:0] = 
0000000000001101010110 + 
1111111111101110111111 = 
{0_1111111111111100010101} < 0
rem[21] = 0000000000001101010110
q = 0000000000000001011000

stage[22]:
force_q_to_zero[22] = ~&(D[31:23]) | ~|(D[22:0]) = 0
{cout[22], sum[22]} = {rem[21], X[9]} + D[22:0] = 
00000000000011010101100 + 
11111111111101110111111 = 
{1_00000000000001001101011} >= 0
rem[22] = 00000000000001001101011
q = 00000000000000010110001

stage[23]:
force_q_to_zero[23] = ~&(D[31:24]) | ~|(D[23:0]) = 0
{cout[23], sum[23]} = {rem[22], X[8]} + D[23:0] = 
000000000000010011010111 + 
111111111111101110111111 = 
{1_000000000000000010010110} >= 0
rem[23] = 000000000000000010010110
q = 000000000000000101100011

stage[24]:
force_q_to_zero[24] = ~&(D[31:25]) | ~|(D[24:0]) = 0
{cout[24], sum[24]} = {rem[23], X[7]} + D[24:0] = 
0000000000000000100101100 + 
1111111111111101110111111 = 
{0_1111111111111110011101011} < 0
rem[24] = 0000000000000000100101100
q = 0000000000000001011000110

stage[25]:
force_q_to_zero[25] = ~&(D[31:26]) | ~|(D[25:0]) = 0
{cout[25], sum[25]} = {rem[24], X[6]} + D[25:0] = 
00000000000000001001011001 + 
11111111111111101110111111 = 
{0_11111111111111111000011000} < 0
rem[25] = 00000000000000001001011001
q = 00000000000000010110001100

stage[26]:
force_q_to_zero[26] = ~&(D[31:27]) | ~|(D[26:0]) = 0
{cout[26], sum[26]} = {rem[25], X[5]} + D[26:0] = 
000000000000000010010110010 + 
111111111111111101110111111 = 
{1_000000000000000000001110001} >= 0
rem[26] = 000000000000000000001110001
q = 000000000000000101100011001

stage[27]:
force_q_to_zero[27] = ~&(D[31:28]) | ~|(D[27:0]) = 0
{cout[27], sum[27]} = {rem[26], X[4]} + D[27:0] = 
0000000000000000000011100010 + 
1111111111111111101110111111 = 
{0_1111111111111111110010100001} < 0
rem[27] = 0000000000000000000011100010
q = 0000000000000001011000110010

stage[28]:
force_q_to_zero[28] = ~&(D[31:29]) | ~|(D[28:0]) = 0
{cout[28], sum[28]} = {rem[27], X[3]} + D[28:0] = 
00000000000000000000111000100 + 
11111111111111111101110111111 = 
{0_11111111111111111110110000011} < 0
rem[28] = 00000000000000000000111000100
q = 00000000000000010110001100100

stage[29]:
force_q_to_zero[29] = ~&(D[31:30]) | ~|(D[29:0]) = 0
{cout[29], sum[29]} = {rem[28], X[2]} + D[29:0] = 
000000000000000000001110001001 + 
111111111111111111101110111111 = 
{0_111111111111111111111101001000} < 0
rem[29] = 000000000000000000001110001001
q = 000000000000000101100011001000

stage[30]:
force_q_to_zero[30] = ~&(D[31:31]) | ~|(D[30:0]) = 0
{cout[30], sum[30]} = {rem[29], X[1]} + D[30:0] = 
0000000000000000000011100010010 + 
1111111111111111111101110111111 = 
{1_0000000000000000000001011010001} >= 0
rem[30] = 0000000000000000000001011010001
q = 0000000000000001011000110010001

stage[31]:
force_q_to_zero[31] = 0
{cout[31], sum[31]} = {rem[30], X[0]} + D[31:0] = 
00000000000000000000010110100011 + 
11111111111111111111101110111111 = 
{1_00000000000000000000000101100010} >= 0
rem[31] = 00000000000000000000000101100010
q = 00000000000000010110001100100011

rem_sign_adj = -rem[31] = 11111111111111111111111010011110

// ---------------------------------------------------------------------------------------------------------------------------------------
由上面的计算过程可知, stage[i](暂时忽略i = 0)需要使用"(i + 1)-bit"的FA来得到q/rem.
设i为整数, 则对于stage[i]和stage[i+1]来说，可以将它们使用的FA都看成"(i + 2)-bit"的(多出来的1-bit宽度正常来说会被EDA优化掉), 即:
for(i = 0; i < 32; i = i + 2)
	Use "(i + 2)-bit" FA for calculation.

在基本的Radix-2 Restoring算法中, 以stage[14, 15]为例:
stage[14]:
temp_rem[14] = {rem[13], X[17]} + (divisor_sign ? D[14:0] : (~D[14:0] + 1'b1))
rem[14] = (temp_rem[14] < 0) ? {rem[13], X[17]} : temp_rem[14];
q[14] = (temp_rem[14] < 0) ? 1'b0 : 1'b1;

stage[15]:
temp_rem[15] = {rem[14], X[16]} + (divisor_sign ? D[15:0] : (~D[15:0] + 1'b1))
rem[15] = (temp_rem[15] < 0) ? {rem[14], X[16]} : temp_rem[15];
q[15] = (temp_rem[15] < 0) ? 1'b0 : 1'b1;

由此可见连续2个"q/rem"的计算是串联的，为了减小延迟，可以并行地计算"q[15, 14]/rem[15, 14]", 对于stage[15], 使用2个FA并行计算"q[14] = 0"和"q[14] = 1"的情况下
temp_rem[15]的值, 即:

temp_rem[15].prev_q_0 = {rem[13], X[17:16]} + (divisor_sign ? D[15:0] : (~D[15:0] + 1'b1));
temp_rem[15].prev_q_1 = {{rem[13], X[17]} + (divisor_sign ? D[14:0] : (~D[14:0] + 1'b1)), X[16]} + (divisor_sign ? D[15:0] : (~D[15:0] + 1'b1));
问题在于计算"temp_rem[15].prev_q_1"的时候，理论上要先做1个3-2 CSA再做1个FA, 这样会导致每2个stage都会引入1个3-2 CSA的延迟.
为了简化描述，将{rem[i], X[30-m]} + (divisor_sign ? D[i+1:0] : (~D[i+1:0] + 1'b1))写为:
{rem[i], X[30-m]} - D[i+1:0]
于是有:
temp_rem[15].prev_q_1 = {({rem[13], X[17]} - D[14:0]), X[16]} - D[15:0] = 
{rem[13], X[17], X[16]} - ({D[14:0], 1'b0} + D[15:0]) = 
{rem[13], X[17:16]} - (3D)[15:0]





3D[(WIDTH + 2)-1:0] = (2D)[(WIDTH + 1)-1:0] + D[WIDTH-1:0] = 
 111111111111111111111011101111110 + 
 111111111111111111111101110111111 = 
1111111111111111111111001100111101
// ---------------------------------------------------------------------------------------------------------------------------------------
写出比较通用的表达式.

for(i = 0; i < WIDTH; i++) begin
	// 边界处的i可能不满足下面的表达式, 暂时忽略
	if(i是偶数) begin
		if(D > 0)
			force_q_to_zero[i] = |(D[(WIDTH-1):(i+1)]);
		else
			// When D < 0, D[WIDTH-1] = 1
			force_q_to_zero[i] = ~&(D[(WIDTH-2):(i+1)]) | ~|(D[i:0]);
		end
	else begin
		if(D > 0) begin
			force_q_to_zero[i].prev_q_0 = |(D[(WIDTH-1):(i+1)]);
			force_q_to_zero[i].prev_q_1 = |(3D[(WIDTH+1):(i+1)]);
		end
		else begin
			// When D < 0, D[WIDTH-1] = 1
			force_q_to_zero[i].prev_q_0 = ~&(D[(WIDTH-2):(i+1)]) | ~|(D[i:0]);
			// When D < 0, 3D[WIDTH+1] = 1
			force_q_to_zero[i].prev_q_1 = ~&(3D[(WIDTH):(i+1)]) | ~|(3D[i:0]);
		end
	end
end




// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
radix-4有符号除法的计算过程:
// ---------------------------------------------------------------------------------------------------------------------------------------
D[WIDTH-1:0] = 11111111111111111111101110111111
abs(X) = 00000101111001101011100101000101
(3D) = 1111111111111111111111001100111101

// ---------------------------
stage[0]:
force_q_to_zero[0] = ~&(D[31:1]) | ~|(D[0:0]) = 1 -> rem[0] = X[31] = 0
q = 0

stage[1]:
force_q_to_zero[1].prev_q_0 = ~&(D[31:2]) | ~|(D[1:0]) = 1
force_q_to_zero[1].prev_q_1 = ~&(3D[32:2]) | ~|(3D[1:0]) = 1

{cout[1].prev_q_0, sum[1].prev_q_0} = {X[31:30]} + D[1:0] = 
00 + 
11 = 
{0_11} < 0
temp_rem[1].prev_q_0 = 00, q[1].prev_q_0 = 0

{cout[1].prev_q_1, sum[1].prev_q_1} = {X[31:30]} + (3D)[1:0] = 
00 + 
01 = 
{0_01} < 0
temp_rem[1].prev_q_1 = 00, q[1].prev_q_1 = 0

q[0] = 0 -> q[1] = q[1].prev_q_0 = 0
q = 00
rem[1] = 00
// ---------------------------
// ---------------------------
stage[2]:
force_q_to_zero[2] = ~&(D[31:3]) | ~|(D[2:0]) = 1
{cout[2], sum[2]} = {rem[1], X[29]} + D[2:0] = 
000 + 
111 = 
{0_111} < 0
rem[2] = 000
q = 000

stage[3]:
force_q_to_zero[3].prev_q_0 = ~&(D[31:4]) | ~|(D[3:0]) = 1
force_q_to_zero[3].prev_q_1 = ~&(3D[32:4]) | ~|(3D[3:0]) = 1

{cout[3].prev_q_0, sum[3].prev_q_0} = {rem[1], X[29:28]} + D[3:0] = 
0000 + 
1111 = 
{0_1111} < 0
temp_rem[3].prev_q_0 = 0000, q[3].prev_q_0 = 0

{cout[3].prev_q_1, sum[3].prev_q_1} = {rem[1], X[29:28]} + (3D)[3:0] = 
0000 + 
1101 = 
{0_1101} < 0
temp_rem[3].prev_q_1 = 0000, q[3].prev_q_1 = 0

q[2] = 0 -> q[3] = q[3].prev_q_0 = 0
q = 0000
rem[3] = 0000
// ---------------------------
// ---------------------------
stage[4]:
force_q_to_zero[4] = ~&(D[31:5]) | ~|(D[4:0]) = 1
{cout[4], sum[4]} = {rem[3], X[27]} + D[4:0] = 
00000 + 
11111 = 
{0_11111} < 0
rem[4] = 00000
q = 00000

stage[5]:
force_q_to_zero[5].prev_q_0 = ~&(D[31:6]) | ~|(D[5:0]) = 1
force_q_to_zero[5].prev_q_1 = ~&(3D[32:6]) | ~|(3D[5:0]) = 1

{cout[5].prev_q_0, sum[5].prev_q_0} = {rem[3], X[27:26]} + D[5:0] = 
000001 + 
111111 = 
{1_000000} >= 0
temp_rem[5].prev_q_0 = 000001, q[5].prev_q_0 = 0

{cout[5].prev_q_1, sum[5].prev_q_1} = {rem[3], X[27:26]} + (3D)[5:0] = 
000001 + 
111101 = 
{0_111110} < 0
temp_rem[5].prev_q_1 = 000001, q[5].prev_q_1 = 0

q[4] = 0 -> q[5] = q[5].prev_q_0 = 0
q = 000000
rem[5] = 000001
// ---------------------------
// ---------------------------
stage[6]:
force_q_to_zero[6] = ~&(D[31:7]) | ~|(D[6:0]) = 1
{cout[6], sum[6]} = {rem[5], X[25]} + D[6:0] = 
0000010 + 
0111111 = 
{0_1000001} < 0
rem[6] = 0000010
q = 0000000

stage[7]:
force_q_to_zero[7].prev_q_0 = ~&(D[31:8]) | ~|(D[7:0]) = 1
force_q_to_zero[7].prev_q_1 = ~&(3D[32:8]) | ~|(3D[7:0]) = 1

{cout[7].prev_q_0, sum[7].prev_q_0} = {rem[5], X[25:24]} + D[7:0] = 
00000101 + 
10111111 = 
{0_11000100} < 0
temp_rem[7].prev_q_0 = 00000101, q[7].prev_q_0 = 0

{cout[7].prev_q_1, sum[7].prev_q_1} = {rem[5], X[25:24]} + (3D)[7:0] = 
00000101 + 
00111101 = 
{0_01000010} < 0
temp_rem[7].prev_q_1 = 00000101, q[7].prev_q_1 = 0

q[6] = 0 -> q[7] = q[7].prev_q_0 = 0
q = 00000000
rem[7] = 00000101
// ---------------------------
// ---------------------------
stage[8]:
force_q_to_zero[8] = ~&(D[31:9]) | ~|(D[8:0]) = 1
{cout[8], sum[8]} = {rem[7], X[23]} + D[8:0] = 
000001011 + 
110111111 = 
{0_111001010} < 0
rem[8] = 000001011
q = 000000000

stage[9]:
force_q_to_zero[9].prev_q_0 = ~&(D[31:10]) | ~|(D[9:0]) = 1
force_q_to_zero[9].prev_q_1 = ~&(3D[32:10]) | ~|(3D[9:0]) = 1

{cout[9].prev_q_0, sum[9].prev_q_0} = {rem[7], X[23:22]} + D[9:0] = 
0000010111 + 
1110111111 = 
{0_1111010110} < 0
temp_rem[9].prev_q_0 = 0000010111, q[9].prev_q_0 = 0

{cout[9].prev_q_1, sum[9].prev_q_1} = {rem[7], X[23:22]} + (3D)[9:0] = 
0000010111 + 
1100111101 = 
{0_1101010100} < 0
temp_rem[9].prev_q_1 = 0000010111, q[9].prev_q_1 = 0

q[8] = 0 -> q[9] = q[9].prev_q_0 = 0
q = 0000000000
rem[9] = 0000010111
// ---------------------------
// ---------------------------
stage[10]:
force_q_to_zero[10] = ~&(D[31:11]) | ~|(D[10:0]) = 0
{cout[10], sum[10]} = {rem[9], X[21]} + D[10:0] = 
00000101111 + 
01110111111 = 
{0_01111101110} < 0
rem[10] = 00000101111
q = 00000000000

stage[11]:
force_q_to_zero[11].prev_q_0 = ~&(D[31:12]) | ~|(D[11:0]) = 0
force_q_to_zero[11].prev_q_1 = ~&(3D[32:12]) | ~|(3D[11:0]) = 0

{cout[11].prev_q_0, sum[11].prev_q_0} = {rem[9], X[21:20]} + D[11:0] = 
000001011110 + 
101110111111 = 
{0_110000011101} < 0
temp_rem[11].prev_q_0 = 000001011110, q[11].prev_q_0 = 0

{cout[11].prev_q_1, sum[11].prev_q_1} = {rem[9], X[21:20]} + (3D)[11:0] = 
000001011110 + 
001100111101 = 
{0_001110011011} < 0
temp_rem[11].prev_q_1 = 000001011110, q[11].prev_q_1 = 0

q[10] = 0 -> q[9] = q[9].prev_q_0 = 0
q = 000000000000
rem[11] = 000001011110
// ---------------------------
// ---------------------------
stage[12]:
force_q_to_zero[12] = ~&(D[31:13]) | ~|(D[12:0]) = 0
{cout[12], sum[12]} = {rem[11], X[19]} + D[12:0] = 
0000010111100 + 
1101110111111 = 
{0_1110001111011} < 0
rem[12] = 0000010111100
q = 0000000000000

stage[13]:
force_q_to_zero[13].prev_q_0 = ~&(D[31:14]) | ~|(D[13:0]) = 0
force_q_to_zero[13].prev_q_1 = ~&(3D[32:14]) | ~|(3D[13:0]) = 0

{cout[13].prev_q_0, sum[13].prev_q_0} = {rem[11], X[19:18]} + D[13:0] = 
00000101111001 + 
11101110111111 = 
{0_11110100111000} < 0
temp_rem[13].prev_q_0 = 00000101111001, q[13].prev_q_0 = 0

{cout[13].prev_q_1, sum[13].prev_q_1} = {rem[11], X[19:18]} + (3D)[13:0] = 
00000101111001 + 
11001100111101 = 
{0_11010010110110} < 0
temp_rem[13].prev_q_1 = 00000101111001, q[13].prev_q_1 = 0

q[12] = 0 -> q[13] = q[13].prev_q_0 = 0
q = 00000000000000
rem[13] = 00000101111001
// ---------------------------
// ---------------------------
stage[14]:
force_q_to_zero[14] = ~&(D[31:15]) | ~|(D[14:0]) = 0
{cout[14], sum[14]} = {rem[13], X[17]} + D[14:0] = 
000001011110011 + 
111101110111111 = 
{0_111111010110010} < 0
rem[14] = 000001011110011
q = 000000000000000

stage[15]:
force_q_to_zero[15].prev_q_0 = ~&(D[31:16]) | ~|(D[15:0]) = 0
force_q_to_zero[15].prev_q_1 = ~&(3D[32:16]) | ~|(3D[15:0]) = 0

{cout[15].prev_q_0, sum[15].prev_q_0} = {rem[13], X[17:16]} + D[15:0] = 
0000010111100110 + 
1111101110111111 = 
{1_0000000110100101} >= 0
temp_rem[15].prev_q_0 = 0000000110100101, q[15].prev_q_0 = 1

{cout[15].prev_q_1, sum[15].prev_q_1} = {rem[13], X[17:16]} + (3D)[15:0] = 
0000010111100110 + 
1111001100111101 = 
{0_1111100100100011} < 0
temp_rem[15].prev_q_1 = 0000010111100110, q[15].prev_q_1 = 0

q[14] = 0 -> q[15] = q[15].prev_q_0 = 1
q = 0000000000000001
rem[15] = 0000000110100101
// ---------------------------
// ---------------------------
stage[16]:
force_q_to_zero[16] = ~&(D[31:17]) | ~|(D[16:0]) = 0
{cout[16], sum[16]} = {rem[15], X[15]} + D[16:0] = 
00000001101001011 + 
11111101110111111 = 
{0_11111111100001010} < 0
rem[16] = 00000001101001011
q = 00000000000000010

stage[17]:
force_q_to_zero[17].prev_q_0 = ~&(D[31:18]) | ~|(D[17:0]) = 0
force_q_to_zero[17].prev_q_1 = ~&(3D[32:18]) | ~|(3D[17:0]) = 0

{cout[17].prev_q_0, sum[17].prev_q_0} = {rem[15], X[15:14]} + D[17:0] = 
000000011010010110 + 
111111101110111111 = 
{1_000000001001010101} >= 0
temp_rem[17].prev_q_0 = 000000001001010101, q[17].prev_q_0 = 1

{cout[17].prev_q_1, sum[17].prev_q_1} = {rem[15], X[15:14]} + (3D)[17:0] = 
000000011010010110 + 
111111001100111101 = 
{0_111111100111010011} < 0
temp_rem[17].prev_q_1 = 000000011010010110, q[17].prev_q_1 = 0

q[16] = 0 -> q[17] = q[16].prev_q_0 = 1
q = 000000000000000101
rem[17] = 000000001001010101
// ---------------------------
// ---------------------------
stage[18]:
force_q_to_zero[18] = ~&(D[31:19]) | ~|(D[18:0]) = 0
{cout[18], sum[18]} = {rem[17], X[13]} + D[18:0] = 
0000000010010101011 + 
1111111101110111111 = 
{1_0000000000001101010} >= 0
rem[18] = 0000000000001101010
q = 0000000000000001011

stage[19]:
force_q_to_zero[19].prev_q_0 = ~&(D[31:20]) | ~|(D[19:0]) = 0
force_q_to_zero[19].prev_q_1 = ~&(3D[32:20]) | ~|(3D[19:0]) = 0

{cout[19].prev_q_0, sum[19].prev_q_0} = {rem[17], X[13:12]} + D[19:0] = 
00000000000011010101 + 
11111111101110111111 = 
{0_11111111110010010100} < 0
temp_rem[19].prev_q_0 = 00000000000011010101, q[19].prev_q_0 = 0

{cout[19].prev_q_1, sum[19].prev_q_1} = {rem[17], X[13:12]} + (3D)[19:0] = 
00000000000011010101 + 
11111111001100111101 = 
{0_111111110100000100100} < 0
temp_rem[19].prev_q_1 = 00000000000011010101, q[19].prev_q_1 = 0

q[18] = 1 -> q[19] = q[19].prev_q_1 = 0
q = 00000000000000010110
rem[19] = 00000000000011010101
// ---------------------------
// ---------------------------
stage[20]:
force_q_to_zero[20] = ~&(D[31:21]) | ~|(D[20:0]) = 0
{cout[20], sum[20]} = {rem[19], X[11]} + D[20:0] = 
000000000000110101011 + 
111111111101110111111 = 
{0_111111111110101101010} < 0
rem[20] = 000000000000110101011
q = 000000000000000101100

stage[21]:
force_q_to_zero[21].prev_q_0 = ~&(D[31:22]) | ~|(D[21:0]) = 0
force_q_to_zero[21].prev_q_1 = ~&(3D[32:22]) | ~|(3D[21:0]) = 0

{cout[21].prev_q_0, sum[21].prev_q_0} = {rem[19], X[11:10]} + D[21:0] = 
0000000000001101010110 + 
1111111111101110111111 = 
{0_1111111111111100010101} < 0
temp_rem[21].prev_q_0 = 0000000000001101010110, q[21].prev_q_0 = 0

{cout[21].prev_q_1, sum[21].prev_q_1} = {rem[19], X[11:10]} + (3D)[21:0] = 
0000000000001101010110 + 
1111111111001100111101 = 
{0_1111111111011010010011} < 0
temp_rem[21].prev_q_1 = 0000000000001101010110, q[21].prev_q_1 = 0

q[20] = 0 -> q[21] = q[21].prev_q_0 = 0
q = 0000000000000001011000
rem[21] = 0000000000001101010110
// ---------------------------
// ---------------------------
stage[22]:
force_q_to_zero[22] = ~&(D[31:23]) | ~|(D[22:0]) = 0
{cout[22], sum[22]} = {rem[21], X[9]} + D[22:0] = 
00000000000011010101100 + 
11111111111101110111111 = 
{1_00000000000001001101011} >= 0
rem[22] = 00000000000001001101011
q = 00000000000000010110001

stage[23]:
force_q_to_zero[23].prev_q_0 = ~&(D[31:24]) | ~|(D[23:0]) = 0
force_q_to_zero[23].prev_q_1 = ~&(3D[32:24]) | ~|(3D[23:0]) = 0

{cout[23].prev_q_0, sum[23].prev_q_0} = {rem[21], X[9:8]} + D[23:0] = 
000000000000110101011001 + 
111111111111101110111111 = 
{1_000000000000100100011000} >= 0
temp_rem[23].prev_q_0 = 000000000000100100011000, q[23].prev_q_0 = 1

{cout[23].prev_q_1, sum[23].prev_q_1} = {rem[21], X[9:8]} + (3D)[23:0] = 
000000000000110101011001 + 
111111111111001100111101 = 
{1_000000000000000010010110} >= 0
temp_rem[23].prev_q_1 = 000000000000000010010110, q[23].prev_q_1 = 1

q[22] = 1 -> q[23] = q[23].prev_q_1 = 1
q = 000000000000000101100011
rem[23] = 000000000000000010010110
// ---------------------------
// ---------------------------
stage[24]:
force_q_to_zero[24] = ~&(D[31:25]) | ~|(D[24:0]) = 0
{cout[24], sum[24]} = {rem[23], X[7]} + D[24:0] = 
0000000000000000100101100 + 
1111111111111101110111111 = 
{0_1111111111111110011101011} < 0
rem[24] = 0000000000000000100101100
q = 0000000000000001011000110

stage[25]:
force_q_to_zero[25].prev_q_0 = ~&(D[31:26]) | ~|(D[25:0]) = 0
force_q_to_zero[25].prev_q_1 = ~&(3D[32:26]) | ~|(3D[25:0]) = 0

{cout[25].prev_q_0, sum[25].prev_q_0} = {rem[23], X[7:6]} + D[25:0] = 
00000000000000001001011001 + 
11111111111111101110111111 = 
{0_11111111111111111000011000} < 0
temp_rem[25].prev_q_0 = 00000000000000001001011001, q[25].prev_q_0 = 0

{cout[25].prev_q_1, sum[25].prev_q_1} = {rem[23], X[7:6]} + (3D)[25:0] = 
00000000000000001001011001 + 
11111111111111001100111101 = 
{0_11111111111111010110010110} < 0
temp_rem[25].prev_q_1 = 00000000000000001001011001, q[25].prev_q_1 = 0

q[24] = 0 -> q[25] = q[25].prev_q_0 = 0
q = 00000000000000010110001100
rem[25] = 00000000000000001001011001
// ---------------------------
// ---------------------------
stage[26]:
force_q_to_zero[26] = ~&(D[31:27]) | ~|(D[26:0]) = 0
{cout[26], sum[26]} = {rem[25], X[5]} + D[26:0] = 
000000000000000010010110010 + 
111111111111111101110111111 = 
{1_000000000000000000001110001} >= 0
rem[26] = 000000000000000000001110001
q = 000000000000000101100011001

stage[27]:
force_q_to_zero[27].prev_q_0 = ~&(D[31:28]) | ~|(D[27:0]) = 0
force_q_to_zero[27].prev_q_1 = ~&(3D[32:28]) | ~|(3D[27:0]) = 0

{cout[27].prev_q_0, sum[27].prev_q_0} = {rem[25], X[5:4]} + D[27:0] = 
0000000000000000100101100100 + 
1111111111111111101110111111 = 
{1_0000000000000000010100100011} >= 0
temp_rem[27].prev_q_0 = 0000000000000000010100100011, q[27].prev_q_0 = 1

{cout[27].prev_q_1, sum[27].prev_q_1} = {rem[25], X[5:4]} + (3D)[27:0] = 
0000000000000000100101100100 + 
1111111111111111001100111101 = 
{0_1111111111111111110010100001} < 0
temp_rem[27].prev_q_1 = 0000000000000000100101100100, q[27].prev_q_1 = 0

q[26] = 1 -> q[27] = q[27].prev_q_1 = 0
q = 0000000000000001011000110010
rem[27] = 0000000000000000000011100010
// ---------------------------
// ---------------------------
stage[28]:
force_q_to_zero[28] = ~&(D[31:29]) | ~|(D[28:0]) = 0
{cout[28], sum[28]} = {rem[27], X[3]} + D[28:0] = 
00000000000000000000111000100 + 
11111111111111111101110111111 = 
{0_11111111111111111110110000011} < 0
rem[28] = 00000000000000000000111000100
q = 00000000000000010110001100100

stage[29]:
force_q_to_zero[29].prev_q_0 = ~&(D[31:30]) | ~|(D[29:0]) = 0
force_q_to_zero[29].prev_q_1 = ~&(3D[32:30]) | ~|(3D[29:0]) = 0

{cout[29].prev_q_0, sum[29].prev_q_0} = {rem[27], X[3:2]} + D[29:0] = 
000000000000000000001110001001 + 
111111111111111111101110111111 = 
{0_111111111111111111111101001000} < 0
temp_rem[29].prev_q_0 = 000000000000000000001110001001, q[29].prev_q_0 = 0

{cout[29].prev_q_1, sum[29].prev_q_1} = {rem[27], X[3:2]} + (3D)[29:0] = 
000000000000000000001110001001 + 
111111111111111111001100111101 = 
{0_111111111111111111011011000110} < 0
temp_rem[29].prev_q_1 = 000000000000000000001110001001, q[29].prev_q_1 = 0

q[28] = 0 -> q[29] = q[28].prev_q_0 = 0
q = 000000000000000101100011001000
rem[29] = 000000000000000000001110001001
// ---------------------------
// ---------------------------
stage[30]:
对于signed_number来说其实不用检测D[31]的值, 如果其是0说明"divisor_is_zero".
force_q_to_zero[30] = ~|(D[30:0]) = 0
{cout[30], sum[30]} = {rem[29], X[1]} + D[30:0] = 
0000000000000000000011100010010 + 
1111111111111111111101110111111 = 
{1_0000000000000000000001011010001} >= 0
rem[30] = 0000000000000000000001011010001
q = 0000000000000001011000110010001

D[WIDTH-1:0] = 11111111111111111111101110111111
abs(X) = 00000101111001101011100101000101
(3D) = 1111111111111111111111001100111101
stage[31]:
force_q_to_zero[31].prev_q_0 = 0
force_q_to_zero[31].prev_q_1 = ~&(3D[32:32]) | ~|(3D[31:0]) = 0

{cout[31].prev_q_0, sum[31].prev_q_0} = {rem[29], X[1:0]} + D[31:0] = 
00000000000000000000111000100101 + 
11111111111111111111101110111111 = 
{1_00000000000000000000100111100100} >= 0
temp_rem[31].prev_q_0 = 00000000000000000000100111100100, q[31].prev_q_0 = 1

{cout[31].prev_q_1, sum[31].prev_q_1} = {rem[29], X[1:0]} + (3D)[31:0] = 
00000000000000000000111000100101 + 
11111111111111111111001100111101 = 
{1_00000000000000000000000101100010} >= 0
temp_rem[31].prev_q_1 = 00000000000000000000000101100010, q[31].prev_q_1 = 1

q[30] = 1 -> q[31] = q[31].prev_q_1 = 1
q = 00000000000000010110001100100011
rem[31] = 00000000000000000000000101100010

rem_sign_adj = -rem[31] = 11111111111111111111111010011110
// ---------------------------





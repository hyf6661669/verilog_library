接"test_1.sv", 此处探究的内容:
将1个或多个"Radix-4"串联起来形成"High-Radix"除法器时，应该如何操作才能得到正确的余数。
对于Radix-N来说, 将Dividend变换到区间"[1/2, 1)"上之后, 需要再向右移:
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N));
N =  4 -> r_shift_num = 1 - ((CLZ_DIFF + 1) % 2);
N =  8 -> r_shift_num = 2 - ((CLZ_DIFF + 1) % 3);
N = 16 -> r_shift_num = 3 - ((CLZ_DIFF + 1) % 4);
N = 32 -> r_shift_num = 4 - ((CLZ_DIFF + 1) % 5);
N = 64 -> r_shift_num = 6 - ((CLZ_DIFF + 1) % 6);
这样最后一次"Radix-N"迭代计算出的"(log2(N))-bit"的商刚好是Q[0 +: log2(N)].
按照上述方法, 做WIDTH-bit整数除法时, 需要用(WIDTH + 1 + 2 + log2(N) - 1) = (WIDTH + 2 + log2(N))来表示w[i].
WIDTH = 32.
假设现在将2个Radix-4串联起来形成Radix-16算法, 即:
N = 16;
(WIDTH + 2 + log2(N)) = 38;

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000000001111111001010100011 = 520867
D[WIDTH-1:0] = 00000000000000000000001011110001 = 753
Q[WIDTH-1:0] = X / D = 691 = 00000000000000000000001010110011
REM[WIDTH-1:0] = 520867 - 753 * 691 = 544 = 00000000000000000000001000100000

CLZ_X = 13
CLZ_D = 22
CLZ_DIFF = CLZ_D - CLZ_X = 9
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (10 % 4) = 1;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(11 / 4) = 3;
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_0111111100101010001100000000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	  = 0_1011110001000000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -17 = 110_1111
m[+0] = - 6 = 111_1001
m[+1] = + 6 = 000_0110
m[+2] = +17 = 001_0001

+ D = 000_1011110001000000000000000000000000000
+2D = 001_0111100010000000000000000000000000000
- D = 111_0100001111000000000000000000000000000
-2D = 110_1000011110000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 1_1100101111000000000000000000000000000 < 0
// 最后一次迭代的商
q_pos = 0100_0000_0100
q_neg = 0001_0101_0000
q_calculated_pre[WIDTH-1:0] = 001010110100
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 001010110011
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
11001011110000000000000000000000 + 10111100010000000000000000000000 = 
10001000000000000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
10001000000000000000000000000000 >> 22 = 
00000000000000000000001000100000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_0001111111001010100011000000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_0111111100101010001100000000000000000
(4 * w[0])_trunc_3_4 = 000_0111, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_0111111100101010001100000000000000000 + 
111_0100001111000000000000000000000000000 = 
111_1100001011101010001100000000000000000 -> 
w[1] = 1_1100001011101010001100000000000000000
4 * w[1] = 111_0000101110101000110000000000000000000
(4 * w[1])_trunc_3_4 = 111_0000, "belongs to [m[-1], m[0])" -> q[2] = -1
q_pos = 0100
q_neg = 0001

// 第2次大迭代
ITER[1]:
4 * w[1] + (-q[2] * D) = 
111_0000101110101000110000000000000000000 + 
000_1011110001000000000000000000000000000 = 
111_1100011111101000110000000000000000000 -> 
w[2] = 1_1100011111101000110000000000000000000
4 * w[2] = 111_0001111110100011000000000000000000000
(4 * w[2])_trunc_3_4 = 111_0001, "belongs to [m[-1], m[0])" -> q[3] = -1
q_pos = 0100_00
q_neg = 0001_01

ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_0001111110100011000000000000000000000 + 
000_1011110001000000000000000000000000000 = 
111_1101101111100011000000000000000000000 -> 
w[3] = 1_1101101111100011000000000000000000000
4 * w[3] = 111_0110111110001100000000000000000000000
(4 * w[3])_trunc_3_4 = 111_0110, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0100_0000
q_neg = 0001_0101

// 第3次大迭代
ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_0110111110001100000000000000000000000 + 
000_1011110001000000000000000000000000000 = 
000_0010101111001100000000000000000000000 -> 
w[4] = 0_0010101111001100000000000000000000000
4 * w[4] = 000_1010111100110000000000000000000000000
(4 * w[4])_trunc_3_4 = 000_1010, "belongs to [m[1], m[2])" -> q[5] = +1
q_pos = 0100_0000_01
q_neg = 0001_0101_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
000_1010111100110000000000000000000000000 + 
111_0100001111000000000000000000000000000 = 
111_1111001011110000000000000000000000000 -> 
w[5] = 1_1111001011110000000000000000000000000
4 * w[5] = 111_1100101111000000000000000000000000000
(4 * w[5])_trunc_3_4 = 111_1100, "belongs to [m[0], m[1])" -> q[6] = 0
q_pos = 0100_0000_0100
q_neg = 0001_0101_0000

// 第4次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
111_1100101111000000000000000000000000000 + 
000_0000000000000000000000000000000000000 = 
111_1100101111000000000000000000000000000 -> 
w[6] = 1_1100101111000000000000000000000000000
4 * w[6] = 111_0010111100000000000000000000000000000
(4 * w[6])_trunc_3_4 = 111_0010, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0100_0000_0100_00
q_neg = 0001_0101_0000_01

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000000011001001001011111010 = 824058
D[WIDTH-1:0] = 00000000000000000000001100000111 = 775
Q[WIDTH-1:0] = X / D = 1063 = 00000000000000000000010000100111
REM[WIDTH-1:0] = 824058 - 775 * 1063 = 233 = 00000000000000000000000011101001

CLZ_X = 12
CLZ_D = 22
CLZ_DIFF = CLZ_D - CLZ_X = 10
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (11 % 4) = 0;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(12 / 4) = 3
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_1100100100101111101000000000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_1100000111000000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -19	= 110_1101
m[+0] = - 6 = 111_1001
m[+1] = + 6 = 000_0110
m[+2] = +19 = 001_0011

+ D = 000_1100000111000000000000000000000000000
+2D = 001_1000001110000000000000000000000000000
- D = 111_0011111001000000000000000000000000000
-2D = 110_0111110010000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6]
w[final] = 0_0011101001000000000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0100_0100_0000
q_neg = 0000_0001_1001
q_calculated_pre[WIDTH-1:0] = 010000100111
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 010000100111
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
00111010010000000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
00111010010000000000000000000000 >> 22 = 
00000000000000000000000011101001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_0011001001001011111010000000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_1100100100101111101000000000000000000
(4 * w[0])_trunc_3_4 = 000_1100, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_1100100100101111101000000000000000000 + 
111_0011111001000000000000000000000000000 = 
000_0000011101101111101000000000000000000 -> 
w[1] = 0_0000011101101111101000000000000000000
4 * w[1] = 000_0001110110111110100000000000000000000
(4 * w[1])_trunc_3_4 = 000_0001, "belongs to [m[0], m[1])" -> q[2] = 0
q_pos = 0100
q_neg = 0000

// 第2次大迭代
ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_0001110110111110100000000000000000000 + 
000_0000000000000000000000000000000000000 = 
000_0001110110111110100000000000000000000 -> 
w[2] = 0_0001110110111110100000000000000000000
4 * w[2] = 000_0111011011111010000000000000000000000
(4 * w[2])_trunc_3_4 = 000_0111, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0100_01
q_neg = 0000_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_0111011011111010000000000000000000000 + 
111_0011111001000000000000000000000000000 = 
111_1011010100111010000000000000000000000 -> 
w[3] = 1_1011010100111010000000000000000000000
4 * w[3] = 110_1101010011101000000000000000000000000
(4 * w[3])_trunc_3_4 = 110_1101, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0100_0100
q_neg = 0000_0001

// 第3次大迭代
ITER[3]:
4 * w[3] + (-q[4] * D) = 
110_1101010011101000000000000000000000000 + 
000_1100000111000000000000000000000000000 = 
111_1001011010101000000000000000000000000 -> 
w[4] = 1_1001011010101000000000000000000000000
4 * w[4] = 110_0101101010100000000000000000000000000
(4 * w[4])_trunc_3_4 = 110_0101, "belongs to [-Inf, m[-1])" -> q[5] = -2
q_pos = 0100_0100_00
q_neg = 0000_0001_10

ITER[4]:
4 * w[4] + (-q[5] * D) = 
110_0101101010100000000000000000000000000 + 
001_1000001110000000000000000000000000000 = 
111_1101111000100000000000000000000000000 -> 
w[5] = 1_1101111000100000000000000000000000000
4 * w[5] = 111_0111100010000000000000000000000000000
(4 * w[5])_trunc_3_4 = 111_0111, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0100_0100_0000
q_neg = 0000_0001_1001

// 第4次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
111_0111100010000000000000000000000000000 + 
000_1100000111000000000000000000000000000 = 
000_0011101001000000000000000000000000000 -> 
w[6] = 0_0011101001000000000000000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000010101010001111001010100011 = 44626595
D[WIDTH-1:0] = 00000000010011001111001011110001 = 5042929
Q[WIDTH-1:0] = X / D = 8 = 00000000000000000000000000001000
REM[WIDTH-1:0] = 44626595 - 5042929 * 8 = 4283163 = 00000000010000010101101100011011

CLZ_X = 6
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 3
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (4 % 4) = 3;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(5 / 4) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_00010101010001111001010100011000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_10011001111001011110001000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -14 = 111_0010
m[+0] = - 4 = 111_1100
m[+1] = + 4	= 000_0100
m[+2] = +14 = 000_1110

+ D = 000_1001100111100101111000100000000000000
+2D = 001_0011001111001011110001000000000000000
- D = 111_0110011000011010000111100000000000000
-2D = 110_1100110000110100001111000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[4];
w[final] = 1_1110100011010000010101000000000000000 < 0
// 最后一次迭代的商
q_pos = 0001_0001
q_neg = 0000_1000
q_calculated_pre[WIDTH-1:0] = 1001
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 1000
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
11101000110100000101010000000000 + 10011001111001011110001000000000
10000010101101100011011000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
10000010101101100011011000000000 >> 9 = 
00000000010000010101101100011011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_0000010101010001111001010100011000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_0001010101000111100101010001100000000
(4 * w[0])_trunc_3_4 = 000_0001, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_0001010101000111100101010001100000000 + 
000_0000000000000000000000000000000000000 = 
000_0001010101000111100101010001100000000 -> 
w[1] = 0_0001010101000111100101010001100000000
4 * w[1] = 000_0101010100011110010101000110000000000
(4 * w[1])_trunc_3_4 = 000_0101, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000

// 第2次大迭代
ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_0101010100011110010101000110000000000 + 
111_0110011000011010000111100000000000000 = 
111_1011101100111000011100100110000000000 -> 
w[2] = 1_1011101100111000011100100110000000000
4 * w[2] = 110_1110110011100001110010011000000000000
(4 * w[2])_trunc_3_4 = 110_1110, "belongs to [-Inf, m[-1])" -> q[3] = -2
q_pos = 0001_00
q_neg = 0000_10

ITER[2]:
4 * w[2] + (-q[3] * D) = 
110_1110110011100001110010011000000000000 + 
001_0011001111001011110001000000000000000 = 
000_0010000010101101100011011000000000000 -> 
w[3] = 0_0010000010101101100011011000000000000
4 * w[3] = 000_1000001010110110001101100000000000000
(4 * w[3])_trunc_3_4 = 000_1000, "belongs to [m[1], m[2])" -> q[4] = +1
q_pos = 0001_0001
q_neg = 0000_1000

// 第3次大迭代
ITER[3]:
4 * w[3] + (-q[4] * D) = 
000_1000001010110110001101100000000000000 + 
111_0110011000011010000111100000000000000 = 
111_1110100011010000010101000000000000000 -> 
w[4] = 1_1110100011010000010101000000000000000

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000111011100000001110100101 = 15598501
D[WIDTH-1:0] = 00000000000000000000000010111011 = 187
Q[WIDTH-1:0] = X / D = 83414 = 00000000000000010100010111010110
REM[WIDTH-1:0] = 44626595 - 187 * 83414 = 83 = 00000000000000000000000001010011

CLZ_X = 8
CLZ_D = 24
CLZ_DIFF = CLZ_D - CLZ_X = 16
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 3 - (17 % 4) = 2;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(18 / 4) = 5
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_0011101110000000111010010100000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_1011101100000000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -17 = 110_1111
m[+0] = - 6 = 111_1010
m[+1] = + 6	= 000_0110
m[+2] = +17 = 000_1110

+ D = 000_1011101100000000000000000000000000000
+2D = 001_0111011000000000000000000000000000000
- D = 111_0100010100000000000000000000000000000
-2D = 110_1000101000000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[10];
w[final] = 0_0101001100000000000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0001_0100_1000_0001_1000
q_neg = 0000_0000_0010_0100_0010
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 00010100010111010110
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 00010100010111010110
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
01010011000000000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
01010011000000000000000000000000 >> 24 = 
00000000000000000000000001010011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_0000111011100000001110100101000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_0011101110000000111010010100000000000
(4 * w[0])_trunc_3_4 = 000_0011, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_0011101110000000111010010100000000000 + 
000_0000000000000000000000000000000000000 = 
000_0011101110000000111010010100000000000 -> 
w[1] = 0_0011101110000000111010010100000000000
4 * w[1] = 000_1110111000000011101001010000000000000
(4 * w[1])_trunc_3_4 = 000_1110, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000

// 第2次大迭代
ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_1110111000000011101001010000000000000 + 
111_0100010100000000000000000000000000000 = 
000_0011001100000011101001010000000000000 -> 
w[2] = 0_0011001100000011101001010000000000000
4 * w[2] = 000_1100110000001110100101000000000000000
(4 * w[2])_trunc_3_4 = 000_1100, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0001_01
q_neg = 0000_00

ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_1100110000001110100101000000000000000 + 
111_0100010100000000000000000000000000000 = 
000_0001000100001110100101000000000000000 -> 
w[3] = 0_0001000100001110100101000000000000000
4 * w[3] = 000_0100010000111010010100000000000000000
(4 * w[3])_trunc_3_4 = 000_0100, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0001_0100
q_neg = 0000_0000

// 第3次大迭代
ITER[3]:
4 * w[3] + (-q[4] * D) = 
000_0100010000111010010100000000000000000 + 
000_0000000000000000000000000000000000000 = 
000_0100010000111010010100000000000000000 -> 
w[4] = 0_0100010000111010010100000000000000000
4 * w[4] = 001_0001000011101001010000000000000000000
(4 * w[4])_trunc_3_4 = 001_0001, "belongs to [m[2], +Inf)" -> q[5] = +2
q_pos = 0001_0100_10
q_neg = 0000_0000_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
001_0001000011101001010000000000000000000 + 
110_1000101000000000000000000000000000000 = 
111_1001101011101001010000000000000000000 -> 
w[5] = 1_1001101011101001010000000000000000000
4 * w[5] = 110_0110101110100101000000000000000000000
(4 * w[5])_trunc_3_4 = 110_0110, "belongs to [-Inf, m[-1])" -> q[6] = -2
q_pos = 0001_0100_1000
q_neg = 0000_0000_0010

// 第4次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
110_0110101110100101000000000000000000000 + 
001_0111011000000000000000000000000000000 = 
111_1110000110100101000000000000000000000 -> 
w[6] = 1_1110000110100101000000000000000000000
4 * w[6] = 111_1000011010010100000000000000000000000
(4 * w[6])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0001_0100_1000_00
q_neg = 0000_0000_0010_01

ITER[6]:
4 * w[6] + (-q[7] * D) = 
111_1000011010010100000000000000000000000 + 
000_1011101100000000000000000000000000000 = 
000_0100000110010100000000000000000000000 -> 
w[7] = 0_0100000110010100000000000000000000000
4 * w[7] = 001_0000011001010000000000000000000000000
(4 * w[7])_trunc_3_4 = 001_0000, "belongs to [m[1], m[2])" -> q[8] = +1
q_pos = 0001_0100_1000_0001
q_neg = 0000_0000_0010_0100

// 第5次大迭代
ITER[7]:
4 * w[7] + (-q[8] * D) = 
001_0000011001010000000000000000000000000 + 
111_0100010100000000000000000000000000000 = 
000_0100101101010000000000000000000000000 -> 
w[8] = 0_0100101101010000000000000000000000000
4 * w[8] = 001_0010110101000000000000000000000000000
(4 * w[8])_trunc_3_4 = 001_0010, "belongs to [m[2], +Inf)" -> q[9] = +2
q_pos = 0001_0100_1000_0001_10
q_neg = 0000_0000_0010_0100_00

ITER[8]:
4 * w[8] + (-q[9] * D) = 
001_0010110101000000000000000000000000000 + 
110_1000101000000000000000000000000000000 = 
111_1011011101000000000000000000000000000 -> 
w[9] = 1_1011011101000000000000000000000000000
4 * w[9] = 110_1101110100000000000000000000000000000
(4 * w[9])_trunc_3_4 = 110_1101, "belongs to [-Inf, m[-1])" -> q[10] = -2
q_pos = 0001_0100_1000_0001_1000
q_neg = 0000_0000_0010_0100_0010

// 第6次大迭代
ITER[9]:
4 * w[9] + (-q[10] * D) = 
110_1101110100000000000000000000000000000 + 
001_0111011000000000000000000000000000000 = 
000_0101001100000000000000000000000000000 -> 
w[10] = 0_0101001100000000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
现在将3个Radix-4串联起来形成Radix-64算法, 即:
N = 64;
(WIDTH + 2 + log2(N)) = 40;

这里有个麻烦的地方, 即log2(64) = 6, 6不是2的幂次, 因此, 对被除数进行规格化操作中的右移步骤中, 右移的位数计算有一定难度。
将CLZ_D = 31 = 1_11111视为特殊情况(这种特殊情况可以通过检查CLZ_D的值是否为全1来获得), 记:
TEMP[5-1:0] = CLZ_DIFF + 1;
则在非特殊(一般)情况下, 必然有:
1 <= TEMP[5-1:0] <= 31
现在的目标是求(TEMP % 6)的值.

按照区间最小值除以8之后向下取整的值，将上述大区间"[1, 31]"划分为以下4个子区间:
1. [ 1,  7]: TEMP[4:3] = 2'd0, TEMP % 6 = TEMP - 0 * 6, OR, TEMP % 6 = TEMP - 1 * 6.
2. [ 8, 15]: TEMP[4:3] = 2'd1, TEMP % 6 = TEMP - 1 * 6, OR, TEMP % 6 = TEMP - 2 * 6.
3. [16, 23]: TEMP[4:3] = 2'd2, TEMP % 6 = TEMP - 2 * 6, OR, TEMP % 6 = TEMP - 3 * 6.
4. [24, 31]: TEMP[4:3] = 2'd3, TEMP % 6 = TEMP - 4 * 6, OR, TEMP % 6 = TEMP - 5 * 6.
因此可以并行计算2个减法:
sub_addend_0[5-1:0] = 
  ({(5){(TEMP[4:3] == 2'd0)}} & 5'd0)
| ({(5){(TEMP[4:3] == 2'd1)}} & 5'd6)
| ({(5){(TEMP[4:3] == 2'd2)}} & 5'd12)
| ({(5){(TEMP[4:3] == 2'd3)}} & 5'd24);
sub_res_0[5-1:0] = TEMP[5-1:0] + ~sub_addend_0[5-1:0] + 5'd1;

sub_addend_1[5-1:0] = 
  ({(5){(TEMP[4:3] == 2'd0)}} & 5'd6)
| ({(5){(TEMP[4:3] == 2'd1)}} & 5'd12)
| ({(5){(TEMP[4:3] == 2'd2)}} & 5'd18)
| ({(5){(TEMP[4:3] == 2'd3)}} & 5'd30);
sub_res_1[6-1:0] = TEMP[5-1:0] + ~sub_addend_1[5-1:0] + 5'd1;

// sub_res_1[5] = 1, 说明"TEMP[5-1:0] >= sub_addend_1[5-1:0]".
TEMP % 6 = sub_res_1[5] ? sub_res_1[3-1:0] : sub_res_0[3-1:0];

以生成TEMP的值开始计算，则得到(TEMP % 6)的延迟包括:
1. 使用TEMP[4:3]生成两个加数, 4选1的Mux.
2. 1个5-bit的全加器.
3. 1个2选1的Mux.

得到(TEMP % 6)之后, 就可以开始右移操作了, 经观察不难发现, 减去6的倍数的操作不会改变(CLZ_DIFF + 1)的LSB的值, 因此在计算(TEMP % 6)的同时也可以执行:
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> (CLZ_DIFF + 1)[0] = 
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> ~CLZ_DIFF[0] = 
得到"r_shift_num = TEMP % 6"之后, 再执行:
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num[2:1];

或者，也可以并行计算两种情况下的右移操作, 即:
Dividend_0 = Dividend >> sub_res_0[2:0];
Dividend_1 = Dividend >> sub_res_1[2:0];
Dividend = sub_res_1[5] ? Dividend_1 : Dividend_0;
对于全加器来说, 结果的LSB肯定比MSB先生成, 因此一般来说算出(sub_res_1[5])的时候"Dividend_0/Dividend_1"的值也得到了....


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000000001111111001010100011 = 520867
D[WIDTH-1:0] = 00000000000000000110000000111111 = 24639
Q[WIDTH-1:0] = X / D = 21 = 00000000000000000000000000010101
REM[WIDTH-1:0] = 520867 - 24639 * 21 = 3448 = 00000000000000000000110101111000

CLZ_X = 13
CLZ_D = 17
CLZ_DIFF = CLZ_D - CLZ_X = 4
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (5 % 6) = 0;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(6 / 6) = 1
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_111111100101010001100000000000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_110000000111111000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -19	= 110_1101
m[+0] = - 6 = 111_1001
m[+1] = + 6 = 000_0110
m[+2] = +19 = 001_0011

+ D = 000_110000000111111000000000000000000000000
+2D = 001_100000001111110000000000000000000000000
- D = 111_001111111000001000000000000000000000000
-2D = 110_011111110000010000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[3];
w[final] = 0_000110101111000000000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0101_01
q_neg = 0000_00
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 010101
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 010101
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
00011010111100000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
00011010111100000000000000000000 >> 17 = 
00000000000000000000110101111000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_001111111001010100011000000000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_111111100101010001100000000000000000000
(4 * w[0])_trunc_3_4 = 000_1111, "belongs to [m[1], m[2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_111111100101010001100000000000000000000 + 
111_001111111000001000000000000000000000000 = 
000_001111011101011001100000000000000000000 -> 
w[1] = 0_001111011101011001100000000000000000000
4 * w[1] = 000_111101110101100110000000000000000000000
(4 * w[1])_trunc_3_4 = 000_1111, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 0101
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_111101110101100110000000000000000000000 + 
111_001111111000001000000000000000000000000 = 
000_001101101101101110000000000000000000000 -> 
w[2] = 0_001101101101101110000000000000000000000
4 * w[2] = 000_110110110110111000000000000000000000000
(4 * w[2])_trunc_3_4 = 000_1101, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0101_01
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_110110110110111000000000000000000000000 + 
111_001111111000001000000000000000000000000 = 
000_000110101111000000000000000000000000000 -> 
w[3] = 0_000110101111000000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000101101100011111011111000 = 11943672
D[WIDTH-1:0] = 00000000000000000101111110100011 = 24483
Q[WIDTH-1:0] = X / D = 487 = 00000000000000000000000111100111
REM[WIDTH-1:0] = 11943672 - 24483 * 487 = 20451 = 00000000000000000100111111100011

CLZ_X = 8
CLZ_D = 17
CLZ_DIFF = CLZ_D - CLZ_X = 9
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (10 % 6) = 1;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(11 / 6) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_010110110001111101111100000000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_101111110100011000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -17 = 110_1111
m[+0] = - 6 = 111_1001
m[+1] = + 6 = 000_0110
m[+2] = +17 = 001_0001

+ D = 000_101111110100011000000000000000000000000
+2D = 001_011111101000110000000000000000000000000
- D = 111_010000001011101000000000000000000000000
-2D = 110_100000010111010000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 1_111000001000000000000000000000000000000 < 0
// 最后一次迭代的商
q_pos = 0010_0000_1000
q_neg = 0000_0010_0000
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 000111101000
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 000111100111
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
11100000100000000000000000000000 + 10111111010001100000000000000000 = 
10011111110001100000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
10011111110001100000000000000000 >> 17 = 
00000000000000000100111111100011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_000101101100011111011111000000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_010110110001111101111100000000000000000
(4 * w[0])_trunc_3_4 = 000_0101, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_010110110001111101111100000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_010110110001111101111100000000000000000 -> 
w[1] = 0_010110110001111101111100000000000000000
4 * w[1] = 001_011011000111110111110000000000000000000
(4 * w[1])_trunc_3_4 = 001_0110, "belongs to [m[2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
001_011011000111110111110000000000000000000 + 
110_100000010111010000000000000000000000000 = 
111_111011011111000111110000000000000000000 -> 
w[2] = 1_111011011111000111110000000000000000000
4 * w[2] = 111_101101111100011111000000000000000000000
(4 * w[2])_trunc_3_4 = 111_1011, "belongs to [m[0], m[1])" -> q[3] = 0
q_pos = 0010_00
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
111_101101111100011111000000000000000000000 + 
000_000000000000000000000000000000000000000 = 
111_101101111100011111000000000000000000000 -> 
w[3] = 1_101101111100011111000000000000000000000
4 * w[3] = 110_110111110001111100000000000000000000000
(4 * w[3])_trunc_3_4 = 110_1101, "belongs to [-Inf, m[-1])" -> q[4] = -2
q_pos = 0010_0000
q_neg = 0000_0010

ITER[3]:
4 * w[3] + (-q[4] * D) = 
110_110111110001111100000000000000000000000 + 
001_011111101000110000000000000000000000000 = 
000_010111011010101100000000000000000000000 -> 
w[4] = 0_010111011010101100000000000000000000000
4 * w[4] = 001_011101101010110000000000000000000000000
(4 * w[4])_trunc_3_4 = 001_0111, "belongs to [m[2], +Inf)" -> q[5] = +2
q_pos = 0010_0000_10
q_neg = 0000_0010_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
001_011101101010110000000000000000000000000 + 
110_100000010111010000000000000000000000000 = 
111_111110000010000000000000000000000000000 -> 
w[5] = 1_111110000010000000000000000000000000000
4 * w[5] = 111_111000001000000000000000000000000000000
(4 * w[5])_trunc_3_4 = 111_1110, "belongs to [m[0], m[1])" -> q[6] = 0
q_pos = 0010_0000_1000
q_neg = 0000_0010_0000

// 第3次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
111_111000001000000000000000000000000000000 + 
000_000000000000000000000000000000000000000 = 
111_111000001000000000000000000000000000000 -> 
w[6] = 1_111000001000000000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000011101100011111011111011 = 7749371
D[WIDTH-1:0] = 00000000000000000101111110100011 = 24483
Q[WIDTH-1:0] = X / D = 316 = 00000000000000000000000100111100
REM[WIDTH-1:0] = 7749371 - 24483 * 316 = 12743 = 00000000000000000011000111000111

CLZ_X = 9
CLZ_D = 17
CLZ_DIFF = CLZ_D - CLZ_X = 8
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (9 % 6) = 2;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(10 / 6) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_001110110001111101111101100000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_101111110100011000000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -17 = 110_1111
m[+0] = - 6 = 111_1001
m[+1] = + 6 = 000_0110
m[+2] = +17 = 001_0001

+ D = 000_101111110100011000000000000000000000000
+2D = 001_011111101000110000000000000000000000000
- D = 111_010000001011101000000000000000000000000
-2D = 110_100000010111010000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 1_101001000100100000000000000000000000000 < 0
// 最后一次迭代的商
q_pos = 0001_0100_0001
q_neg = 0000_0000_0100
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 000100111101
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 000100111100
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
10100100010010000000000000000000 + 10111111010001100000000000000000 = 
01100011100011100000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
01100011100011100000000000000000 >> 17 = 
00000000000000000011000111000111 = REM[WIDTH-1:0]
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_000011101100011111011111011000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_001110110001111101111101100000000000000
(4 * w[0])_trunc_3_4 = 000_0011, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_001110110001111101111101100000000000000 + 
000_000000000000000000000000000000000000000 = 
000_001110110001111101111101100000000000000 -> 
w[1] = 0_001110110001111101111101100000000000000
4 * w[1] = 000_111011000111110111110110000000000000000
(4 * w[1])_trunc_3_4 = 000_1110, "belongs to [m[1], m[2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_111011000111110111110110000000000000000 + 
111_010000001011101000000000000000000000000 = 
000_001011010011011111110110000000000000000 -> 
w[2] = 0_001011010011011111110110000000000000000
4 * w[2] = 000_101101001101111111011000000000000000000
(4 * w[2])_trunc_3_4 = 000_1011, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0001_01
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_101101001101111111011000000000000000000 + 
111_010000001011101000000000000000000000000 = 
111_111101011001100111011000000000000000000 -> 
w[3] = 1_111101011001100111011000000000000000000
4 * w[3] = 111_110101100110011101100000000000000000000
(4 * w[3])_trunc_3_4 = 111_1101, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0001_0100
q_neg = 0000_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_110101100110011101100000000000000000000 + 
000_000000000000000000000000000000000000000 = 
111_110101100110011101100000000000000000000 -> 
w[4] = 1_110101100110011101100000000000000000000
4 * w[4] = 111_010110011001110110000000000000000000000
(4 * w[4])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[5] = -1
q_pos = 0001_0100_00
q_neg = 0000_0000_01

ITER[4]:
4 * w[4] + (-q[5] * D) = 
111_010110011001110110000000000000000000000 + 
000_101111110100011000000000000000000000000 = 
000_000110001110001110000000000000000000000 -> 
w[5] = 0_000110001110001110000000000000000000000
4 * w[5] = 000_011000111000111000000000000000000000000
(4 * w[5])_trunc_3_4 = 000_0110, "belongs to [m[1], m[2])" -> q[6] = +1
q_pos = 0001_0100_0001
q_neg = 0000_0000_0100

// 第3次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
000_011000111000111000000000000000000000000 + 
111_010000001011101000000000000000000000000 = 
111_101001000100100000000000000000000000000 -> 
w[6] = 1_101001000100100000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000011101100011111011111011 = 7749371
D[WIDTH-1:0] = 00000000000000001111000110100011 = 61859
Q[WIDTH-1:0] = X / D = 125 = 00000000000000000000000001111101
REM[WIDTH-1:0] = 7749371 - 61859 * 125 = 16996 = 00000000000000000100001001100100

CLZ_X = 9
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 7
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (8 % 6) = 3;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(9 / 6) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_000111011000111110111110110000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_111100011010001100000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -24 = 110_1000
m[+0] = - 8 = 111_1000
m[+1] = + 8 = 000_1000
m[+2] = +24 = 001_1000

+ D = 000_111100011010001100000000000000000000000
+2D = 001_111000110100011000000000000000000000000
- D = 111_000011100101110100000000000000000000000
-2D = 110_000111001011101000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 0_010000100110010000000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0000_1000_0001
q_neg = 0000_0000_0100
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 01111101
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 01111101
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
01000010011001000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
01000010011001000000000000000000 >> 16 = 
00000000000000000100001001100100 = REM[WIDTH-1:0]
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_000001110110001111101111101100000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_000111011000111110111110110000000000000
(4 * w[0])_trunc_3_4 = 000_0001, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_000111011000111110111110110000000000000 + 
000_000000000000000000000000000000000000000 = 
000_000111011000111110111110110000000000000 -> 
w[1] = 0_000111011000111110111110110000000000000
4 * w[1] = 000_011101100011111011111011000000000000000
(4 * w[1])_trunc_3_4 = 000_0111, "belongs to [m[0], m[1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_011101100011111011111011000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_011101100011111011111011000000000000000 -> 
w[2] = 0_011101100011111011111011000000000000000
4 * w[2] = 001_110110001111101111101100000000000000000
(4 * w[2])_trunc_3_4 = 001_1101, "belongs to [m[2], +Inf)" -> q[3] = +2
q_pos = 0000_10
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
001_110110001111101111101100000000000000000 + 
110_000111001011101000000000000000000000000 = 
111_111101011011010111101100000000000000000 -> 
w[3] = 1_111101011011010111101100000000000000000
4 * w[3] = 111_110101101101011110110000000000000000000
(4 * w[3])_trunc_3_4 = 111_1101, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0000_1000
q_neg = 0000_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_110101101101011110110000000000000000000 + 
110_000111001011101000000000000000000000000 = 
111_110101101101011110110000000000000000000 -> 
w[4] = 1_110101101101011110110000000000000000000
4 * w[4] = 111_010110110101111011000000000000000000000
(4 * w[4])_trunc_3_4 = 111_0101, "belongs to [m[-1], m[0])" -> q[5] = -1
q_pos = 0000_1000_00
q_neg = 0000_0000_01

ITER[4]:
4 * w[4] + (-q[5] * D) = 
111_010110110101111011000000000000000000000 + 
000_111100011010001100000000000000000000000 = 
000_010011010000000111000000000000000000000 -> 
w[5] = 0_010011010000000111000000000000000000000
4 * w[5] = 001_001101000000011100000000000000000000000
(4 * w[5])_trunc_3_4 = 001_0011, "belongs to [m[1], m[2])" -> q[6] = +1
q_pos = 0000_1000_0001
q_neg = 0000_0000_0100

// 第3次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
001_001101000000011100000000000000000000000 + 
111_000011100101110100000000000000000000000 = 
000_010000100110010000000000000000000000000 -> 
w[6] = 0_010000100110010000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000001101100011111011111011 = 3555067
D[WIDTH-1:0] = 00000000000000001111000110100011 = 61859
Q[WIDTH-1:0] = X / D = 57 = 00000000000000000000000000111001
REM[WIDTH-1:0] = 3555067 - 61859 * 57 = 29104 = 00000000000000000111000110110000

CLZ_X = 10
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 6
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (7 % 6) = 4;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(8 / 6) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_000011011000111110111110110000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_111100011010001100000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -24 = 110_1000
m[+0] = - 8 = 111_1000
m[+1] = + 8 = 000_1000
m[+2] = +24 = 001_1000

+ D = 000_111100011010001100000000000000000000000
+2D = 001_111000110100011000000000000000000000000
- D = 111_000011100101110100000000000000000000000
-2D = 110_000111001011101000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 0_011100011011000000000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0000_0100_0001
q_neg = 0000_0000_1000
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 00111001
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 00111001
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
01110001101100000000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
01110001101100000000000000000000 >> 16 = 
00000000000000000111000110110000 = REM[WIDTH-1:0]
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_000000110110001111101111101100000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_000011011000111110111110110000000000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_000011011000111110111110110000000000000 + 
000_000000000000000000000000000000000000000 = 
000_000011011000111110111110110000000000000 -> 
w[1] = 0_000011011000111110111110110000000000000
4 * w[1] = 000_001101100011111011111011000000000000000
(4 * w[1])_trunc_3_4 = 000_0011, "belongs to [m[0], m[1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_001101100011111011111011000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_001101100011111011111011000000000000000 -> 
w[2] = 0_001101100011111011111011000000000000000
4 * w[2] = 000_110110001111101111101100000000000000000
(4 * w[2])_trunc_3_4 = 000_1101, "belongs to [m[1], m[2])" -> q[3] = +1
q_pos = 0000_01
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_110110001111101111101100000000000000000 + 
111_000011100101110100000000000000000000000 = 
111_111001110101100011101100000000000000000 -> 
w[3] = 1_111001110101100011101100000000000000000
4 * w[3] = 111_100111010110001110110000000000000000000
(4 * w[3])_trunc_3_4 = 111_1001, "belongs to [m[0], m[1])" -> q[4] = 0
q_pos = 0000_0100
q_neg = 0000_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
111_100111010110001110110000000000000000000 + 
000_000000000000000000000000000000000000000 = 
111_100111010110001110110000000000000000000 -> 
w[4] = 1_100111010110001110110000000000000000000
4 * w[4] = 110_011101011000111011000000000000000000000
(4 * w[4])_trunc_3_4 = 110_0111, "belongs to [-Inf, m[-1])" -> q[5] = -2
q_pos = 0000_0100_00
q_neg = 0000_0000_10

ITER[4]:
4 * w[4] + (-q[5] * D) = 
110_011101011000111011000000000000000000000 + 
001_111000110100011000000000000000000000000 = 
000_010110001101010011000000000000000000000 -> 
w[5] = 0_010110001101010011000000000000000000000
4 * w[5] = 001_011000110101001100000000000000000000000
(4 * w[5])_trunc_3_4 = 001_0110, "belongs to [m[1], m[2])" -> q[6] = +1
q_pos = 0000_0100_0001
q_neg = 0000_0000_1000

// 第3次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
001_011000110101001100000000000000000000000 + 
111_000011100101110100000000000000000000000 = 
000_011100011011000000000000000000000000000 -> 
w[6] = 0_011100011011000000000000000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 00000000000111111111111111111000 = 2097144
D[WIDTH-1:0] = 00000000000000001111000110100011 = 61859
Q[WIDTH-1:0] = X / D = 33 = 00000000000000000000000000100001
REM[WIDTH-1:0] = 2097144 - 61859 * 33 = 55797 = 00000000000000001101100111110101

CLZ_X = 11
CLZ_D = 16
CLZ_DIFF = CLZ_D - CLZ_X = 5
被除数规格化操作步骤:
1. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, X[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}}, 小数点在"Dividend[MSB], Dividend[MSB-1]"之间.
2. r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % 6) = 5 - (6 % 6) = 5;
3. Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] >> r_shift_num;
除数规格化操作步骤:
1. Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = {1'b0, D[WIDTH-1:0] << CLZ_X, {(2 + log2(N) - 1){1'b0}}};
需要迭代的次数:
iter_num = ceil((CLZ_DIFF + 1 + 1) / log2(N)) = ceil(7 / 6) = 2
Dividend[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_000001111111111111111110000000000000000
Divisor[(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] 	= 0_111100011010001100000000000000000000000
根据Divisor的值, 可得选择常数:
m[-1] = -24 = 110_1000
m[+0] = - 8 = 111_1000
m[+1] = + 8 = 000_1000
m[+2] = +24 = 001_1000

+ D = 000_111100011010001100000000000000000000000
+2D = 001_111000110100011000000000000000000000000
- D = 111_000011100101110100000000000000000000000
-2D = 110_000111001011101000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6];
w[final] = 0_110110011111010100000000000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0000_0010_00_01
q_neg = 0000_0000_00_00
q_calculated_pre[WIDTH-1:0] = q_pos - q_neg = 00100001
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] - (w[final] < 0) = 00100001
remainder_calculated_pre[WIDTH-1:0] = w[final][(2 + log2(N) - 1) +: WIDTH] + ((w[final] < 0) ? Divisor[(2 + log2(N) - 1) +: WIDTH] : {(WIDTH){1'b0}}) = 
11011001111101010000000000000000
remainder_calculated[WIDTH-1:0] = remainder_calculated_pre[WIDTH-1:0] >> CLZ_D = 
11011001111101010000000000000000 >> 16 = 
00000000000000001101100111110101 = REM[WIDTH-1:0]
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w[0][(WIDTH + 1 + 2 + (log2(N) - 1))-1:0] = Dividend / 4 = 0_000000011111111111111111100000000000000
q[0] = 0

// 第1次大迭代
4 * w[0] = 000_000001111111111111111110000000000000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
4 * w[0] + (-q[1] * D) = 
000_000001111111111111111110000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_000001111111111111111110000000000000000 -> 
w[1] = 0_000001111111111111111110000000000000000
4 * w[1] = 000_000111111111111111111000000000000000000
(4 * w[1])_trunc_3_4 = 000_0001, "belongs to [m[0], m[1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
4 * w[1] + (-q[2] * D) = 
000_000111111111111111111000000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_000111111111111111111000000000000000000 -> 
w[2] = 0_000111111111111111111000000000000000000
4 * w[2] = 000_011111111111111111100000000000000000000
(4 * w[2])_trunc_3_4 = 000_0111, "belongs to [m[0], m[1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00

// 第2次大迭代
ITER[2]:
4 * w[2] + (-q[3] * D) = 
000_011111111111111111100000000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_011111111111111111100000000000000000000 -> 
w[3] = 0_011111111111111111100000000000000000000
4 * w[3] = 001_111111111111111110000000000000000000000
(4 * w[3])_trunc_3_4 = 001_1111, "belongs to [m[2], +Inf)" -> q[4] = +2
q_pos = 0000_0010
q_neg = 0000_0000

ITER[3]:
4 * w[3] + (-q[4] * D) = 
001_111111111111111110000000000000000000000 + 
110_000111001011101000000000000000000000000 = 
000_000111001011100110000000000000000000000 -> 
w[4] = 0_000111001011100110000000000000000000000
4 * w[4] = 000_011100101110011000000000000000000000000
(4 * w[4])_trunc_3_4 = 000_0111, "belongs to [m[0], m[1])" -> q[5] = 0
q_pos = 0000_0010_00
q_neg = 0000_0000_00

ITER[4]:
4 * w[4] + (-q[5] * D) = 
000_011100101110011000000000000000000000000 + 
000_000000000000000000000000000000000000000 = 
000_011100101110011000000000000000000000000 -> 
w[5] = 0_011100101110011000000000000000000000000
4 * w[5] = 001_110010111001100000000000000000000000000
(4 * w[5])_trunc_3_4 = 001_1100, "belongs to [m[1], m[2])" -> q[6] = +1
q_pos = 0000_0010_00_01
q_neg = 0000_0000_00_00

// 第3次大迭代
ITER[5]:
4 * w[5] + (-q[6] * D) = 
001_110010111001100000000000000000000000000 + 
111_000011100101110100000000000000000000000 = 
000_110110011111010100000000000000000000000 -> 
w[6] = 0_110110011111010100000000000000000000000









算是人工验证完毕了吧...


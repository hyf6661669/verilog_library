测试使用Divisor取反后的值来进行迭代，是否还能得到正确的结果
WIDTH = 28;


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110100001110011100100011 = 13690659
D[WIDTH-1:0] = 0000000000001010000000000000 = 40960
Q[WIDTH-1:0] = X / D = 334 = 0000000000000000000101001110
REM[WIDTH-1:0] = 13690659 - 40960 * 334 = 10019 = 0000000000000010011100100011

CLZ_X = 4
CLZ_D = 12
CLZ_DIFF = CLZ_D - CLZ_X = 8
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (9 % 2) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(10 / 2) = 5;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 1101000011100111001000110000
Divisor[WIDTH-1:0] 		= 1010000000000000000000000000

+ D = 0_1010000000000000000000000000000
+2D = 1_0100000000000000000000000000000
- D = 1_0110000000000000000000000000000
-2D = 0_1100000000000000000000000000000
~ D = 1_0101111111111111111111111111111
~2D = 0_1011111111111111111111111111111

4 * (+ D) = 010_1000000000000000000000000000000
4 * (+2D) = 101_0000000000000000000000000000000
4 * (~ D) = 101_0111111111111111111111111111100
4 * (~2D) = 010_1111111111111111111111111111100

根据D的值, 可得选择常数:
m[-1] = -16 = 111_0000
m[ 0] = - 6 = 111_1010
m[+1] = + 6 = 000_0110
m[+2] = +16 = 001_0000

-m[-1]_reduced_2_5 = 01_00000
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 11_00000

// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[5];
w[5] = 4 * w[4] - q[5] * D = 
1_0110011100100011000000000000000 + 
0_1100000000000000000000000000000 = 
0_0010011100100011000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0101_0100_10
q_neg = 0000_0001_00
corr(q_pos - q_neg) = 000101001110

w[final]_reduced >> CLZ_D = 0010011100100011000000000000 >> 12 = 
0000000000000010011100100011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// REM是负数
REM = -10019 = 1111111111111101100011011101
w_sum[4] = 0_1010010000110111001111111111000
w_carry[4] = 1_1011010110010001100000000001000
4 * w_sum[4] = 0_1001000011011100111111111100000
4 * w_carry[4] = 0_1101011001000110000000000100000
-q[5] * D = -2D = 0_1100000000000000000000000000000


(~0_1001000011011100111111111100000 + 1) + (~0_1101011001000110000000000100000 + 1) + (~0_1100000000000000000000000000000 + 1) = 
(1_0110111100100011000000000100000 + 1_0010100110111001111111111100000 + 1_0100000000000000000000000000000)_reduced = 
1_1101100011011101000000000000

(1_1101100011011101000000000000 / (2 ^ CLZ_D))_reduced = 
1111111111111101100011011101
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


初始化:
w_sum[0] 	= 0_0011010000111001110010001100000
w_carry[0] 	= 0_0000000000000000000000000000000
w[0] = 0_0011010000111001110010001100000
(4 * w[0])_trunc_3_4 = 000_1101, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00


ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
1_1000111100011000110111001111111
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_1010000111001110010001100000001
w[1] = 4 * w[0] - q[1] * D = 
0_1101000011100111001000110000000 + 
1_0110000000000000000000000000000 = 
0_0011000011100111001000110000000
(4 * w[1])_trunc_3_4 = 000_1100, "belongs to [m[+1], m[+2])" -> q[2] = +1
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
110_0011 + 010_1000 = 000_1011, "belongs to [m[+1], m[+2])" -> q[2] = +1


// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_01000 + 00_00000 + 01_00000 = 00_01000
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_0100 + 000_0000 + 000_0110 = 011_1010
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_0100 + 000_0000 + 111_1010 = 010_1110
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_01000 + 00_00000 + 11_00000 = 10_01000


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (00_01000 + 01_01111)_reduced_2_4 = 
(01_10111)_reduced_2_4 = 01_1011 >= 0, don't care.
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (011_1010 + 101_0111)_reduced_3_3 = 
(001_0001)_reduced_3_3 = 001_000 >= 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (010_1110 + 101_0111)_reduced_3_3 = 
(11_10111)_reduced_3_3 = 11_1011 < 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_01000 + 01_01111)_reduced_2_4 = 
(11_00000)_reduced_2_4 = 11_0000 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0101
q_neg = 0000


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
1_1110010010100101100101000000111
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_0011111011110110111101111111001
w[2] = 4 * w[1] - q[2] * D = 
0_1100001110011100100011000000000 + 
1_0110000000000000000000000000000 = 
0_0010001110011100100011000000000
(4 * w[2])_trunc_3_4 = 000_1000, "belongs to [m[+1], m[+2])" -> q[3] = +1
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
111_1001 + 000_1111 = 000_1000, "belongs to [m[+1], m[+2])" -> q[3] = +1


// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_11110 + 10_00011 + 01_00000 = 00_00001
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
000_1111 + 010_0001 + 000_0110 = 011_0110
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
000_1111 + 010_0001 + 111_1010 = 010_1010
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_11110 + 10_00011 + 11_00000 = 10_00001


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (00_00001 + 01_01111)_reduced_2_4 = 
(01_10000)_reduced_2_4 = 01_1000 >= 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (011_0110 + 101_0111)_reduced_3_3 = 
(000_1101)_reduced_3_3 = 000_110 >= 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (010_1010 + 101_0111)_reduced_3_3 = 
(000_0001)_reduced_3_3 = 000_000 >= 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (10_00001 + 01_01111)_reduced_2_4 = 
(11_10000)_reduced_2_4 = 11_1000 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[3] = +1
q_pos = 0101_01
q_neg = 0000_00


ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_0011011010110010011100000000111
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
1_1011011110111111101111111111001
w[3] = 4 * w[2] - q[3] * D = 
0_1000111001110010001100000000000 + 
1_0110000000000000000000000000000 = 
1_1110111001110010001100000000000
(4 * w[3])_trunc_3_4 = 111_1011, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0101_0100
q_neg = 0000_0000
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_1101 + 110_1101 = 111_1010, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0101_0100
q_neg = 0000_0000

// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_01001 + 11_11101 + 01_00000 = 11_00110
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_0100 + 011_1110 + 000_0110 = 010_1000
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_0100 + 011_1110 + 111_1010 = 001_1100
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_01001 + 11_11101 + 11_00000 = 01_00110


(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (11_00110 + 01_01111)_reduced_2_4 = 
(00_10101)_reduced_2_4 = 00_1010 >= 0
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (010_1000 + 101_0111)_reduced_3_3 = 
(111_1111)_reduced_3_3 = 111_111 < 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (001_1100 + 101_0111)_reduced_3_3 = 
(111_0011)_reduced_3_3 = 111_001 < 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (01_00110 + 01_01111)_reduced_2_4 = 
(10_10101)_reduced_2_4 = 10_1010 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[4] = -1
q_pos = 0101_0100
q_neg = 0000_0001


ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_1010010000110111001111111111000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_1011010110010001100000000001000
w[4] = 4 * w[3] - q[4] * D = 
1_1011100111001000110000000000000 + 
0_1010000000000000000000000000000 = 
0_0101100111001000110000000000000
(4 * w[4])_trunc_3_4 = 001_0110, "belongs to [m[+2], +Inf)" -> q[5] = +2
q_pos = 0101_0100_10
q_neg = 0000_0001_00
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
010_1001 + 110_1101 = 001_0110, "belongs to [m[+2], +Inf)" -> q[5] = +2
q_pos = 0101_0100_10
q_neg = 0000_0001_00

// From the paper:
temp[4][0] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_01101 + 11_01111 + 01_00000 = 11_11100
temp[4][1] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_0110 + 011_0111 + 000_0110 = 111_0011
temp[4][2] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_0110 + 011_0111 + 111_1010 = 110_0111
temp[4][3] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_01101 + 11_01111 + 11_00000 = 01_11100

4 * (+ D) = 00010_10000000000000000000000000000
(temp[4][0] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (11_11100 + 10_10000)_reduced_2_4 = 
(10_01100)_reduced_2_4 = 10_0110 < 0, don't care.
(temp[4][1] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (111_0011 + 010_1000)_reduced_3_3 = 
(001_1011)_reduced_3_3 = 001_101 >= 0
(temp[4][2] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (110_0111 + 010_1000)_reduced_3_3 = 
(000_1111)_reduced_3_3 = 000_111 >= 0
(temp[4][3] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (01_11100 + 10_10000)_reduced_2_4 = 
(00_01100)_reduced_2_4 = 00_0110 >= 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+2], +Inf)" -> q[5] = +2
q_pos = 0101_0100_10
q_neg = 0000_0001_00


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1000010110011111011100111011 = 140113723
D[WIDTH-1:0] = 0000000000000110000001000011 = 24643
Q[WIDTH-1:0] = X / D = 5685 = 0000000000000001011000110101
REM[WIDTH-1:0] = 140113723 - 24643 * 5685 = 18268 = 0000000000000100011101011100

CLZ_X = 0
CLZ_D = 13
CLZ_DIFF = CLZ_D - CLZ_X = 13
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (14 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(15 / 2) = 8;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000010110011111011100111011
Divisor[WIDTH-1:0] 		= 1100000010000110000000000000

+ D = 0_1100000010000110000000000000000
+2D = 1_1000000100001100000000000000000
- D = 1_0011111101111010000000000000000
-2D = 0_0111111011110100000000000000000
~ D = 1_0011111101111001111111111111111
~2D = 0_0111111011110011111111111111111

4 * (+ D) = 011_0000001000011000000000000000000
4 * (+2D) = 110_0000010000110000000000000000000
4 * (~ D) = 100_1111110111100111111111111111100
4 * (~2D) = 001_1111101111001111111111111111100

根据D的值, 可得选择常数:
m[-1] = -18 = 110_1110
m[ 0] = - 6 = 111_1010
m[+1] = + 6 = 000_0110
m[+2] = +18 = 001_0010

-m[-1]_reduced_2_5 = 01_00100
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 10_11100

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8];
w[8] = 4 * w[7] - q[8] * D = 
1_0100111100111110000000000000000 + 
0_0111111011110100000000000000000 = 
1_1100111000110010000000000000000 < 0
// 最后一次迭代的商
q_pos = 0001_1000_0100_0110
q_neg = 0000_0010_0001_0000
corr(q_pos - q_neg) = 0001011000110101

(w[final]_reduced + (+D)) >> CLZ_D = 
(1100111000110010000000000000 + 1100000010000110000000000000) >> 13 = 
1000111010111000000000000000 >> 13 = 
0000000000000100011101011100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// REM是负数
REM = -18268 = 1111111111111011100010100100
w_sum[7] = 1_1011010101101100100000000111111
w_carry[7] = 0_1001111001100010111111111000001
4 * w_sum[7] = 0_1101010110110010000000011111100
4 * w_carry[7] = 0_0111100110001011111111100000100
-q[8] * D = -2D = 0_0111111011110100000000000000000


(~0_1101010110110010000000011111100 + 1) + (~0_0111100110001011111111100000100 + 1) + (~0_0111111011110100000000000000000 + 1) = 
(1_0010101001001101111111100000100 + 1_1000011001110100000000011111100 + 1_1000000100001100000000000000000)_reduced = 
0_0011000111001110000000000000

0_0011000111001110000000000000 + (-D) = 
0_0011000111001110000000000000 + 1_0011111101111010000000000000 = 
1_0111000101001000000000000000

(1_0111000101001000000000000000 / (2 ^ CLZ_D))_reduced = 
1111111111111011100010100100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] 	= 0_0001000010110011111011100111011
w_carry[0] 	= 0_0000000000000000000000000000000
w[0] = 0_0001000010110011111011100111011
(4 * w[0])_trunc_3_4 = 000_0100, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00


ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_0100001011001111101110011101100
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_0000000000000000000000000000000
w[1] = 4 * w[0] - q[1] * D = 
0_0100001011001111101110011101100 + 
0_0000000000000000000000000000000 = 
0_0100001011001111101110011101100
(4 * w[1])_trunc_3_4 = 001_0000, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
001_0000 + 000_0000 = 001_0000, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_00001 + 00_00000 + 01_00100 = 10_00101
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_0000 + 000_0000 + 000_0110 = 001_0110
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_0000 + 000_0000 + 111_1010 = 000_1010
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_00001 + 00_00000 + 10_11100 = 11_11101


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_00101 + 00_00000)_reduced_2_4 = 
(10_00101)_reduced_2_4 = 10_0010 < 0, don't care.
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (001_0110 + 000_0000)_reduced_3_3 = 
(001_0110)_reduced_3_3 = 001_011 >= 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (000_1010 + 000_0000)_reduced_3_3 = 
(000_1010)_reduced_3_3 = 000_1010 >= 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (11_11101 + 00_00000)_reduced_2_4 = 
(11_11101)_reduced_2_4 = 11_1110 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[2] = +1
q_pos = 0001
q_neg = 0000


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_0011010001000111000110001001111
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_0001011001110001110011101100001
w[2] = 4 * w[1] - q[2] * D = 
1_0000101100111110111001110110000 + 
1_0011111101111010000000000000000 = 
0_0100101010111000111001110110000
(4 * w[2])_trunc_3_4 = 001_0010, "belongs to [m[+2], +Inf)" -> q[3] = +2
q_pos = 0001_10
q_neg = 0000_00
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_1101 + 000_0101 = 001_0010, "belongs to [m[+2], +Inf)" -> q[3] = +2
q_pos = 0001_10
q_neg = 0000_00


// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
00_00101 + 00_00000 + 01_00100 = 01_01001
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
100_0010 + 000_0000 + 000_0110 = 100_1000
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
100_0010 + 000_0000 + 111_1010 = 011_1100
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
00_00101 + 00_00000 + 10_11100 = 11_00001


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (01_01001 + 00_11111)_reduced_2_4 = 
(10_01000)_reduced_2_4 = 10_0100 < 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (100_1000 + 100_1111)_reduced_3_3 = 
(001_0111)_reduced_3_3 = 001_011 >= 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (011_1100 + 100_1111)_reduced_3_3 = 
(000_1011)_reduced_3_3 = 000_101 >= 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (11_00001 + 00_11111)_reduced_2_4 = 
(00_00000)_reduced_2_4 = 00_0000 >= 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+2], +Inf)" -> q[3] = +2
q_pos = 0001_10
q_neg = 0000_00


ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_1111011000101000101001101000111
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_1011001110101110111101101111001
w[3] = 4 * w[2] - q[3] * D = 
1_0010101011100011100111011000000 + 
0_0111111011110100000000000000000 = 
1_1010100111010111100111011000000
(4 * w[3])_trunc_3_4 = 110_1010, "belongs to (-Inf, m[-1])" -> q[4] = -2
q_pos = 0001_1000
q_neg = 0000_0010
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
011_1101 + 010_1100 = 101_1001, "belongs to (-Inf, m[-1])" -> q[4] = -2
q_pos = 0001_1000
q_neg = 0000_0010


// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_01000 + 01_01100 + 01_00100 = 01_11000
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_0100 + 001_0110 + 000_0110 = 101_0000
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_0100 + 001_0110 + 111_1010 = 100_0100
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_01000 + 01_01100 + 10_11100 = 11_10000


(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (01_11000 + 01_11111)_reduced_2_4 = 
(11_10111)_reduced_2_4 = 11_1011 < 0
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (101_0000 + 001_1111)_reduced_3_3 = 
(110_1111)_reduced_3_3 = 110_111 < 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (100_0100 + 001_1111)_reduced_3_3 = 
(110_0011)_reduced_3_3 = 110_001 < 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (11_10000 + 01_11111)_reduced_2_4 = 
(01_01111)_reduced_2_4 = 01_0111 >= 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to (-Inf, m[-1])" -> q[4] = -2
q_pos = 0001_1000
q_neg = 0000_0010


ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_1001011100010101010000011111000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_1001000101010101001101000001000
w[4] = 4 * w[3] - q[4] * D = 
0_1010011101011110011101100000000 + 
1_1000000100001100000000000000000 = 
0_0010100001101010011101100000000
(4 * w[4])_trunc_3_4 = 000_1010, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0001_1000_01
q_neg = 0000_0010_00
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
010_0101 + 110_0100 = 000_1001, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0001_1000_01
q_neg = 0000_0010_00


// From the paper:
temp[4][0] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_01100 + 11_00111 + 01_00100 = 11_10111
temp[4][1] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
111_0110 + 011_0011 + 000_0110 = 010_1111
temp[4][2] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
111_0110 + 011_0011 + 111_1010 = 010_0011
temp[4][3] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_01100 + 11_00111 + 10_11100 = 01_01111


(temp[4][0] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (11_10111 + 10_00000)_reduced_2_4 = 
(01_10111)_reduced_2_4 = 01_1011 >= 0, don't care.
(temp[4][1] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (010_1111 + 110_0000)_reduced_3_3 = 
(000_1111)_reduced_3_3 = 000_111 >= 0
(temp[4][2] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (010_0011 + 110_0000)_reduced_3_3 = 
(000_0011)_reduced_3_3 = 000_001 >= 0
(temp[4][3] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (01_01111 + 10_00000)_reduced_2_4 = 
(11_01111)_reduced_2_4 = 11_0111 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0001_1000_01
q_neg = 0000_0010_00


ITER[4]:
w_sum[5] = csa_sum(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
1_0010011001111000001010000111111
w_carry[5] = csa_carry(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
0_1011101010101011101011111000001
w[5] = 4 * w[4] - q[5] * D = 
0_1010000110101001110110000000000 + 
1_0011111101111010000000000000000 = 
1_1110000100100011110110000000000
(4 * w[5])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0001_1000_0100
q_neg = 0000_0010_0001
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
100_1001 + 010_1110 = 111_0111, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0001_1000_0100
q_neg = 0000_0010_0001


// From the paper:
temp[5][0] = ((16 * w_sum[4])_reduced_2_5 + (16 * w_carry[4])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_01110 + 01_00010 + 01_00100 = 11_10100
temp[5][1] = ((16 * w_sum[4])_reduced_3_4 + (16 * w_carry[4])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_0111 + 001_0001 + 000_0110 = 010_1110
temp[5][2] = ((16 * w_sum[4])_reduced_3_4 + (16 * w_carry[4])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_0111 + 001_0001 + 111_1010 = 010_0010
temp[5][3] = ((16 * w_sum[4])_reduced_2_5 + (16 * w_carry[4])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_01110 + 01_00010 + 10_11100 = 01_01100


(temp[5][0] + (-4 * q[5] * D)_reduced_2_5)_reduced_2_4 = (11_10100 + 00_11111)_reduced_2_4 = 
(00_10011)_reduced_2_4 = 00_1001 >= 0
(temp[5][1] + (-4 * q[5] * D)_reduced_3_4)_reduced_3_3 = (010_1110 + 100_1111)_reduced_3_3 = 
(111_1101)_reduced_3_3 = 111_110 < 0
(temp[5][2] + (-4 * q[5] * D)_reduced_3_4)_reduced_3_3 = (010_0010 + 100_1111)_reduced_3_3 = 
(111_0001)_reduced_3_3 = 111_000 < 0
(temp[5][3] + (-4 * q[5] * D)_reduced_2_5)_reduced_2_4 = (01_01100 + 00_11111)_reduced_2_4 = 
(10_01011)_reduced_2_4 = 10_0101 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[6] = -1
q_pos = 0001_1000_0100
q_neg = 0000_0010_0001


ITER[5]:
w_sum[6] = csa_sum(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
0_1011001111001000000111111111000
w_carry[6] = csa_carry(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
1_1001000101001101010000000001000
w[6] = 4 * w[5] - q[6] * D = 
1_1000010010001111011000000000000 + 
0_1100000010000110000000000000000 = 
0_0100010100010101011000000000000
(4 * w[6])_trunc_3_4 = 001_0001, "belongs to [m[+1], m[+2])" -> q[7] = +1
q_pos = 0001_1000_0100_01
q_neg = 0000_0010_0001_00
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
010_1100 + 110_0100 = 001_0000, "belongs to [m[+1], m[+2])" -> q[7] = +1
q_pos = 0001_1000_0100_01
q_neg = 0000_0010_0001_00


// From the paper:
temp[6][0] = ((16 * w_sum[5])_reduced_2_5 + (16 * w_carry[5])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_01100 + 11_10101 + 01_00100 = 11_00101
temp[6][1] = ((16 * w_sum[5])_reduced_3_4 + (16 * w_carry[5])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
010_0110 + 011_1010 + 000_0110 = 110_0110
temp[6][2] = ((16 * w_sum[5])_reduced_3_4 + (16 * w_carry[5])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
010_0110 + 011_1010 + 111_1010 = 101_1010
temp[6][3] = ((16 * w_sum[5])_reduced_2_5 + (16 * w_carry[5])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_01100 + 11_10101 + 10_11100 = 00_11101


(temp[6][0] + (-4 * q[6] * D)_reduced_2_5)_reduced_2_4 = (11_00101 + 11_00000)_reduced_2_4 = 
(10_00101)_reduced_2_4 = 10_0010 < 0, don't care.
(temp[6][1] + (-4 * q[6] * D)_reduced_3_4)_reduced_3_3 = (110_0110 + 011_0000)_reduced_3_3 = 
(001_0110)_reduced_3_3 = 001_011 >= 0
(temp[6][2] + (-4 * q[6] * D)_reduced_3_4)_reduced_3_3 = (101_1010 + 011_0000)_reduced_3_3 = 
(000_1010)_reduced_3_3 = 000_101 >= 0
(temp[6][3] + (-4 * q[6] * D)_reduced_2_5)_reduced_2_4 = (00_11101 + 11_00000)_reduced_2_4 = 
(11_11101)_reduced_2_4 = 11_1110 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[7] = +1
q_pos = 0001_1000_0100_01
q_neg = 0000_0010_0001_00


ITER[6]:
w_sum[7] = csa_sum(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
1_1011010101101100100000000111111
w_carry[7] = csa_carry(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
0_1001111001100010111111111000001
w[7] = 4 * w[6] - q[7] * D = 
1_0001010001010101100000000000000 + 
1_0011111101111010000000000000000 = 
0_0101001111001111100000000000000
(4 * w[7])_trunc_3_4 = 001_0100, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0001_1000_0100_0110
q_neg = 0000_0010_0001_0000
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
110_1101 + 010_0111 = 001_0100, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0001_1000_0100_0110
q_neg = 0000_0010_0001_0000


// From the paper:
temp[7][0] = ((16 * w_sum[6])_reduced_2_5 + (16 * w_carry[6])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_00111 + 01_00010 + 01_00100 = 01_01101
temp[7][1] = ((16 * w_sum[6])_reduced_3_4 + (16 * w_carry[6])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_0011 + 001_0001 + 000_0110 = 100_1010
temp[7][2] = ((16 * w_sum[6])_reduced_3_4 + (16 * w_carry[6])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_0011 + 001_0001 + 111_1010 = 011_1110
temp[7][3] = ((16 * w_sum[6])_reduced_2_5 + (16 * w_carry[6])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_00111 + 01_00010 + 10_11100 = 11_00101

4 * (~ D) = 100_1111110111100111111111111111100
(temp[7][0] + (-4 * q[7] * D)_reduced_2_5)_reduced_2_4 = (01_01101 + 00_11111)_reduced_2_4 = 
(10_01100)_reduced_2_4 = 10_0110 < 0, don't care.
(temp[7][1] + (-4 * q[7] * D)_reduced_3_4)_reduced_3_3 = (100_1010 + 100_1111)_reduced_3_3 = 
(001_1001)_reduced_3_3 = 001_100 >= 0
(temp[7][2] + (-4 * q[7] * D)_reduced_3_4)_reduced_3_3 = (011_1110 + 100_1111)_reduced_3_3 = 
(000_1101)_reduced_3_3 = 000_110 >= 0
(temp[7][3] + (-4 * q[7] * D)_reduced_2_5)_reduced_2_4 = (11_00101 + 00_11111)_reduced_2_4 = 
(00_00100)_reduced_2_4 = 00_0010 >= 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+2], +Inf)" -> q[8] = +2
q_pos = 0001_1000_0100_0110
q_neg = 0000_0010_0001_0000


// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------

WIDTH = 32
1 + WIDTH + 2 + 1 = 36

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 01010000110100001110011100100011 = 1355867939
D[WIDTH-1:0] = 00000000101000000000100000000011 = 10487811
Q[WIDTH-1:0] = X / D = 129 = 00000000000000000000000010000001
REM[WIDTH-1:0] = 1355867939 - 10487811 * 129 = 2940320 = 00000000001011001101110110100000

CLZ_X = 1
CLZ_D = 8
CLZ_DIFF = CLZ_D - CLZ_X = 7
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (8 % 2) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(9 / 2) = 5;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 10100001101000011100111001000110
Divisor[WIDTH-1:0] 		= 10100000000010000000001100000000

+ D = 0_10100000000010000000001100000000000
+2D = 1_01000000000100000000011000000000000
- D = 1_01011111111101111111110100000000000
-2D = 0_10111111111011111111101000000000000
~ D = 1_01011111111101111111110011111111111
~2D = 0_10111111111011111111100111111111111

4 * (+ D) = 010_10000000001000000000110000000000000
4 * (+2D) = 101_00000000010000000001100000000000000
4 * (~ D) = 101_01111111110111111111001111111111100
4 * (~2D) = 010_11111111101111111110011111111111100

根据D的值, 可得选择常数:
m[-1] = -16 = 111_0000
m[ 0] = - 6 = 111_1010
m[+1] = + 6 = 000_0110
m[+2] = +16 = 001_0000

-m[-1]_reduced_2_5 = 01_00000
-m[ 0]_reduced_3_4 = 000_0110
-m[+1]_reduced_3_4 = 111_1010
-m[+2]_reduced_2_5 = 11_00000

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[5];
w[5] = 4 * w[4] - q[5] * D = 
0_11001100111001011010001100000000000 + 
1_01011111111101111111110100000000000 = 
0_00101100110111011010000000000000000 >= 0
// 最后一次迭代的商
q_pos = 0010_0000_01
q_neg = 0000_0000_00
corr(q_pos - q_neg) = 0010000001

w[final]_reduced >> CLZ_D = 00101100110111011010000000000000 >> 8 = 
00000000001011001101110110100000
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] 	= 0_00010100001101000011100111001000110
w_carry[0] 	= 0_00000000000000000000000000000000000
w[0] = 0_00010100001101000011100111001000110
(4 * w[0])_trunc_3_4 = 000_0101, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_01010000110100001110011100100011000
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000000000000000
w[1] = 4 * w[0] - q[1] * D = 
0_01010000110100001110011100100011000 + 
0_00000000000000000000000000000000000 = 
0_01010000110100001110011100100011000
(4 * w[1])_trunc_3_4 = 001_0100, "belongs to [m[+2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_01000 + 00_00000 + 01_00000 = 10_01000
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
001_0100 + 000_0000 + 000_0110 = 001_1010
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
001_0100 + 000_0000 + 111_1010 = 000_1110
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_01000 + 00_00000 + 11_00000 = 00_01000


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_01000 + 00_00000)_reduced_2_4 = 
(10_01000)_reduced_2_4 = 10_0100 < 0, don't care.
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (001_1010 + 000_0000)_reduced_3_3 = 
(001_1010)_reduced_3_3 = 001_101 >= 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (000_1110 + 000_0000)_reduced_3_3 = 
(000_1110)_reduced_3_3 = 000_111 >= 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (00_01000 + 00_00000)_reduced_2_4 = 
(00_01000)_reduced_2_4 = 00_0100 >= 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+2], +Inf)" -> q[2] = +2
q_pos = 0010
q_neg = 0000


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
1_11111100101011000110010101110011111
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_00000110100001110011000100011000001
w[2] = 4 * w[1] - q[2] * D = 
1_01000011010000111001110010001100000 + 
0_10111111111011111111101000000000000 = 
0_00000011001100111001011010001100000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0010_00
q_neg = 0000_00

// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_00001 + 00_00000 + 01_00000 = 10_00001
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
101_0000 + 000_0000 + 000_0110 = 101_0110
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
101_0000 + 000_0000 + 111_1010 = 100_1010
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_00001 + 00_00000 + 11_00000 = 00_00001


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (10_00001 + 10_11111)_reduced_2_4 = 
(01_00000)_reduced_2_4 = 01_0000 >= 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (101_0110 + 010_1111)_reduced_3_3 = 
(000_0101)_reduced_3_3 = 000_010 >= 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (100_1010 + 010_1111)_reduced_3_3 = 
(111_1001)_reduced_3_3 = 111_100 < 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (00_00001 + 10_11111)_reduced_2_4 = 
(11_00000)_reduced_2_4 = 11_0000 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0010_00
q_neg = 0000_00


ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
1_11101000101011010101000110101111000
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_00100100001000010000100010000001000
w[3] = 4 * w[2] - q[3] * D = 
0_00001100110011100101101000110000000 + 
0_00000000000000000000000000000000000 = 
0_00001100110011100101101000110000000
(4 * w[3])_trunc_3_4 = 000_0011, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0010_0000
q_neg = 0000_0000

// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_11001 + 00_01101 + 01_00000 = 01_00110
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
111_1100 + 000_0110 + 000_0110 = 000_1000
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
111_1100 + 000_0110 + 111_1010 = 111_1100
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_11001 + 00_01101 + 11_00000 = 11_00110


(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (01_00110 + 00_00000)_reduced_2_4 = 
(01_00110)_reduced_2_4 = 01_0011 >= 0, don't care.
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (000_1000 + 000_0000)_reduced_3_3 = 
(000_1000)_reduced_3_3 = 000_100 >= 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (111_1100 + 000_0000)_reduced_3_3 = 
(111_1100)_reduced_3_3 = 111_110 < 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (11_00110 + 00_00000)_reduced_2_4 = 
(11_00110)_reduced_2_4 = 11_0011 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0010_0000
q_neg = 0000_0000


ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_00110010001100010110010010111000000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_00000001000010000000010000001000000
w[4] = 4 * w[3] - q[4] * D = 
0_00110011001110010110100011000000000 + 
0_00000000000000000000000000000000000 = 
0_00110011001110010110100011000000000
(4 * w[4])_trunc_3_4 = 000_1100, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0010_0000_01
q_neg = 0000_0000_00

// From the paper:
temp[4][0] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_10001 + 10_01000 + 01_00000 = 01_11001
temp[4][1] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_1000 + 010_0100 + 000_0110 = 001_0010
temp[4][2] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_1000 + 010_0100 + 111_1010 = 000_0110
temp[4][3] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_10001 + 10_01000 + 11_00000 = 11_11001


(temp[4][0] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (01_11001 + 00_00000)_reduced_2_4 = 
(01_11001)_reduced_2_4 = 01_1100 >= 0, don't care.
(temp[4][1] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (001_0010 + 000_0000)_reduced_3_3 = 
(001_0010)_reduced_3_3 = 001_001 >= 0
(temp[4][2] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (000_0110 + 000_0000)_reduced_3_3 = 
(000_0110)_reduced_3_3 = 000_011 >= 0
(temp[4][3] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (11_11001 + 00_00000)_reduced_2_4 = 
(11_11001)_reduced_2_4 = 11_1100 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0010_0000_01
q_neg = 0000_0000_00



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 01110110110100010000011110111001 = 1993410489
D[WIDTH-1:0] = 00000000011110000000000000000000 = 7864320
Q[WIDTH-1:0] = X / D = 253 = 00000000000000000000000011111101
REM[WIDTH-1:0] = 1993410489 - 7864320 * 253 = 3737529 = 00000000001110010000011110111001

CLZ_X = 1
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 8
r_shift_num = log2(N) - 1 - ((CLZ_DIFF + 1) % log2(N)) = 1 - (9 % 2) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 2) / log2(N)) = ceil(10 / 2) = 5;

规格化操作之后:
Dividend[WIDTH-1:0] 	= 11101101101000100000111101110010
Divisor[WIDTH-1:0] 		= 11110000000000000000000000000000

+ D = 0_11110000000000000000000000000000000
+2D = 1_11100000000000000000000000000000000
- D = 1_00010000000000000000000000000000000
-2D = 0_00100000000000000000000000000000000
~ D = 1_00001111111111111111111111111111111
~2D = 0_00011111111111111111111111111111111

4 * (+ D) = 011_11000000000000000000000000000000000
4 * (+2D) = 111_10000000000000000000000000000000000
4 * (~ D) = 100_00111111111111111111111111111111100
4 * (~2D) = 000_01111111111111111111111111111111100

根据D的值, 可得选择常数:
m[-1] = -23 = 110_1001
m[ 0] = - 8 = 111_1000
m[+1] = + 8 = 000_1000
m[+2] = +23 = 001_0111

-m[-1]_reduced_2_5 = 01_01110
-m[ 0]_reduced_3_4 = 000_1000
-m[+1]_reduced_3_4 = 111_1000
-m[+2]_reduced_2_5 = 10_10010

// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[5];
w[5] = 4 * w[4] - q[5] * D = 
1_01100010000011110111001000000000000 + 
1_00010000000000000000000000000000000 = 
0_01110010000011110111001000000000000 >= 0
// 最后一次迭代的商
q_pos = 0100_0000_01
q_neg = 0000_0001_00
corr(q_pos - q_neg) = 11111101

w[final]_reduced >> CLZ_D = 01110010000011110111001000000000 >> 9 = 
00000000001110010000011110111001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w_sum[0] 	= 0_00111011011010001000001111011100100
w_carry[0] 	= 0_00000000000000000000000000000000000
w[0] = 0_00111011011010001000001111011100100
(4 * w[0])_trunc_3_4 = 000_1110, "belongs to [m[+1], m[+2])" -> q[1] = +1
q_pos = 01
q_neg = 00

ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
1_11100010010111011111000010001101111
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_00011011010001000001111011100100001
w[1] = 4 * w[0] - q[1] * D = 
0_11101101101000100000111101110010000 + 
1_00010000000000000000000000000000000 = 
1_11111101101000100000111101110010000
(4 * w[1])_trunc_3_4 = 111_1111, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0100
q_neg = 0000

// From the paper:
temp[1][0] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
11_10110 + 00_00000 + 01_01110 = 01_00100
temp[1][1] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
011_1011 + 000_0000 + 000_1000 = 100_0011
temp[1][2] = ((16 * w_sum[0])_reduced_3_4 + (16 * w_carry[0])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
011_1011 + 000_0000 + 111_1000 = 011_0011
temp[1][3] = ((16 * w_sum[0])_reduced_2_5 + (16 * w_carry[0])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
11_10110 + 00_00000 + 10_10010 = 10_01000


(temp[1][0] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (01_00100 + 00_00111)_reduced_2_4 = 
(11_10011)_reduced_2_4 = 11_1001 < 0, don't care.
(temp[1][1] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (100_0011 + 100_0011)_reduced_3_3 = 
(000_0110)_reduced_3_3 = 000_011 >= 0
(temp[1][2] + (-4 * q[1] * D)_reduced_3_4)_reduced_3_3 = (011_0011 + 100_0011)_reduced_3_3 = 
(111_0110)_reduced_3_3 = 111_011 < 0
(temp[1][3] + (-4 * q[1] * D)_reduced_2_5)_reduced_2_4 = (10_01000 + 00_00111)_reduced_2_4 = 
(10_01111)_reduced_2_4 = 10_0111 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0100
q_neg = 0000


ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
1_11100100011001111011100110100111000
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_00010010001000001000010000100001000
w[2] = 4 * w[1] - q[2] * D = 
1_11110110100010000011110111001000000 + 
0_00000000000000000000000000000000000 = 
1_11110110100010000011110111001000000
(4 * w[2])_trunc_3_4 = 111_1101, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0100_00
q_neg = 0000_00

// From the paper:
temp[2][0] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_00100 + 01_10110 + 01_01110 = 01_01000
temp[2][1] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_0010 + 001_1011 + 000_1000 = 000_0101
temp[2][2] = ((16 * w_sum[1])_reduced_3_4 + (16 * w_carry[1])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_0010 + 001_1011 + 111_1000 = 111_0101
temp[2][3] = ((16 * w_sum[1])_reduced_2_5 + (16 * w_carry[1])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_00100 + 01_10110 + 10_10010 = 10_01100


(temp[2][0] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (01_01000 + 00_00000)_reduced_2_4 = 
(01_01000)_reduced_2_4 = 01_0100 >= 0, don't care.
(temp[2][1] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (000_0101 + 000_0000)_reduced_3_3 = 
(000_0101)_reduced_3_3 = 000_010 >= 0
(temp[2][2] + (-4 * q[2] * D)_reduced_3_4)_reduced_3_3 = (111_0101 + 000_0000)_reduced_3_3 = 
(111_0101)_reduced_3_3 = 111_010 < 0
(temp[2][3] + (-4 * q[2] * D)_reduced_2_5)_reduced_2_4 = (10_01100 + 00_00000)_reduced_2_4 = 
(10_01100)_reduced_2_4 = 10_0110 < 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0100_00
q_neg = 0000_00


ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
1_11011001000111001111011000011000000
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_00000001000001000000000100001000000
w[3] = 4 * w[2] - q[3] * D = 
1_11011010001000001111011100100000000 + 
0_00000000000000000000000000000000000 = 
1_11011010001000001111011100100000000
(4 * w[3])_trunc_3_4 = 111_0110, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0100_0000
q_neg = 0000_0001

// From the paper:
temp[3][0] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
10_01000 + 01_00100 + 01_01110 = 00_11010
temp[3][1] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
110_0100 + 001_0010 + 000_1000 = 111_1110
temp[3][2] = ((16 * w_sum[2])_reduced_3_4 + (16 * w_carry[2])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
110_0100 + 001_0010 + 111_1000 = 110_1110
temp[3][3] = ((16 * w_sum[2])_reduced_2_5 + (16 * w_carry[2])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
10_01000 + 01_00100 + 10_10010 = 01_11110


(temp[3][0] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (00_11010 + 00_00000)_reduced_2_4 = 
(00_11010)_reduced_2_4 = 00_1101 >= 0
(temp[3][1] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (111_1110 + 000_0000)_reduced_3_3 = 
(111_1110)_reduced_3_3 = 111_111 < 0
(temp[3][2] + (-4 * q[3] * D)_reduced_3_4)_reduced_3_3 = (110_1110 + 000_0000)_reduced_3_3 = 
(110_1110)_reduced_3_3 = 110_111 < 0
(temp[3][3] + (-4 * q[3] * D)_reduced_2_5)_reduced_2_4 = (01_11110 + 00_00000)_reduced_2_4 = 
(01_11110)_reduced_2_4 = 01_1111 >= 0, don't care.
根据比较结果(Sign Detection, SD)可得, "belongs to [m[-1], m[0])" -> q[4] = -1
q_pos = 0100_0000
q_neg = 0000_0001


ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
1_11011001000111001111011000011000000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_00000001000001000000000100001000000
w[4] = 4 * w[3] - q[4] * D = 
1_01101000100000111101110010000000000 + 
0_11110000000000000000000000000000000 = 
0_01011000100000111101110010000000000
(4 * w[4])_trunc_3_4 = 001_0110, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0100_0000_01
q_neg = 0000_0001_00

// From the paper:
temp[4][0] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[-1]_reduced_2_5)_reduced_2_5 = 
01_10010 + 00_00010 + 01_01110 = 11_00010
temp[4][1] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[ 0]_reduced_3_4)_reduced_3_4 = 
101_1001 + 000_0001 + 000_1000 = 110_0010
temp[4][2] = ((16 * w_sum[3])_reduced_3_4 + (16 * w_carry[3])_reduced_3_4 + -m[+1]_reduced_3_4)_reduced_3_4 = 
101_1001 + 000_0001 + 111_1000 = 101_0010
temp[4][3] = ((16 * w_sum[3])_reduced_2_5 + (16 * w_carry[3])_reduced_2_5 + -m[+2]_reduced_2_5)_reduced_2_5 = 
01_10010 + 00_00010 + 10_10010 = 00_00110


(temp[4][0] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (11_00010 + 11_11000)_reduced_2_4 = 
(10_11010)_reduced_2_4 = 10_1101 < 0, don't care.
(temp[4][1] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (110_0010 + 011_1100)_reduced_3_3 = 
(001_1110)_reduced_3_3 = 001_111 >= 0
(temp[4][2] + (-4 * q[4] * D)_reduced_3_4)_reduced_3_3 = (101_0010 + 011_1100)_reduced_3_3 = 
(000_1110)_reduced_3_3 = 000_111 >= 0
(temp[4][3] + (-4 * q[4] * D)_reduced_2_5)_reduced_2_4 = (00_00110 + 11_11000)_reduced_2_4 = 
(11_11110)_reduced_2_4 = 11_1111 < 0
根据比较结果(Sign Detection, SD)可得, "belongs to [m[+1], m[+2])" -> q[5] = +1
q_pos = 0100_0000_01
q_neg = 0000_0001_00



+ D = 0_10000000000000000000000000000000000
~ D = 1_01111111111111111111111111111111111
- D = 1_10000000000000000000000000000000000
sum = 0_00010000000000000000000000000000000
cry = 0_00000000000000000000000000000000000

0_01000000000000000000000000000000000
1_01111111111111111111111111111111111

sum_o = 1_00111111111111111111111111111111111
cry_o = 0_10000000000000000000000000000000001


sum = 0_00100000000000000000000000000000000
cry = 0_00000000000000000000000000000000000
+ D = 0_11111111111111111111111111111111000
- D = 1_00000000000000000000000000000001000
~ D = 1_00000000000000000000000000000000111

0_10000000000000000000000000000000000
1_00000000000000000000000000000000111

sum_o = 1_10000000000000000000000000000000111
cry_o = 0_00000000000000000000000000000000001


w = 
0_10000000000000000000000000000000000 + 
1_00000000000000000000000000000001000 = 
1_10000000000000000000000000000001000
测试"WIDTH = 16"时, 使用"WIDTH = 32"的计算模块进行SRT迭代的设计.
这次使用"sum/carry"来进行中间迭代, 测试将位宽扩大之后，最后是否只需要使用16-bit的FA就能算出余数.

// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 16;
ITN = InTerNal
ITN_W = 1 + (2 * WIDTH) = 33;
0_00000000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0001010010010100 = 5268
D[WIDTH-1:0] = 0000001000000011 = 515
Q[WIDTH-1:0] = X / D = 10 = 0000000000001010
REM[WIDTH-1:0] = 5268 - 515 * 10 = 118 = 0000000001110110

CLZ_X = 3
CLZ_D = 6
CLZ_DIFF = CLZ_D - CLZ_X = 3
Normalized_D = 1000000011000000
根据D的值, 可得选择常数:
m[-1] = -13
m[ 0] = - 4
m[+1] = + 4
m[+2] = +12

+ D[ITN_W-1:0] = 0_10000000110000000000000000000000
+2D[ITN_W-1:0] = 1_00000001100000000000000000000000
- D[ITN_W-1:0] = 1_01111111010000000000000000000000
-2D[ITN_W-1:0] = 0_11111110100000000000000000000000
~ D[ITN_W-1:0] = 1_01111111001111111111111111111111
~2D[ITN_W-1:0] = 0_11111110011111111111111111111111

l_shift_num = CLZ_D = 6
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_00000000000000000001010010010100 << 6 = 
0_00000000000001010010010100000000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w_sum[0][ITN_W-1:0] 	= 0_00000000000001010010010100000000
w_carry[0][ITN_W-1:0] 	= 0_00000000000000000000000000000000
w[0] 					= 0_00000000000001010010010100000000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_00000000000101001001010000000000
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_00000000000000000000000000000000
w[1] = w[0] << 2 - q[1] * D = 
0_00000000000101001001010000000000 + 
0_00000000000000000000000000000000 = 
0_00000000000101001001010000000000
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_00000000010100100101000000000000
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_00000000000000000000000000000000
w[2] = w[1] << 2 - q[2] * D = 
0_00000000010100100101000000000000 + 
0_00000000000000000000000000000000 = 
0_00000000010100100101000000000000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00

ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_00000001010010010100000000000000
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_00000000000000000000000000000000
w[3] = w[2] << 2 - q[3] * D = 
0_00000001010010010100000000000000 + 
0_00000000000000000000000000000000 = 
0_00000001010010010100000000000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000

ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_00000101001001010000000000000000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_00000000000000000000000000000000
w[4] = w[3] << 2 - q[4] * D = 
0_00000101001001010000000000000000 + 
0_00000000000000000000000000000000 = 
0_00000101001001010000000000000000
(4 * w[4])_trunc_3_4 = 000_0001, "belongs to [m[0], m[+1])" -> q[5] = 0
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00

ITER[4]:
w_sum[5] = csa_sum(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
0_00010100100101000000000000000000
w_carry[5] = csa_carry(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
0_00000000000000000000000000000000
w[5] = w[4] << 2 - q[5] * D = 
0_00010100100101000000000000000000 + 
0_00000000000000000000000000000000 = 
0_00010100100101000000000000000000
(4 * w[5])_trunc_3_4 = 000_0101, "belongs to [m[+1], m[+2])" -> q[6] = +1
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
000_0101 + 000_0000 = 000_0101, "belongs to [m[+1], m[+2])" -> q[6] = +1
q_pos = 0000_0000_0001
q_neg = 0000_0000_0000

ITER[5]:
w_sum[6] = csa_sum(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
1_00101101011011111111111111111111
w_carry[6] = csa_carry(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
0_10100100001000000000000000000001
w[6] = w[5] << 2 - q[6] * D = 
0_01010010010100000000000000000000 + 
1_01111111010000000000000000000000 = 
1_11010001100100000000000000000000
(4 * w[6])_trunc_3_4 = 111_0100, "belongs to [m[-1], m[0])" -> q[7] = -1
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
100_1011 + 010_1001 = 111_0100, "belongs to [m[-1], m[0])" -> q[7] = -1
q_pos = 0000_0000_0001_00
q_neg = 0000_0000_0000_01

ITER[6]:
w_sum[7] = csa_sum(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
0_10100101111111111111111111111000
w_carry[7] = csa_carry(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
1_00100001000000000000000000001000
w[7] = w[6] << 2 - q[7] * D = 
1_01000110010000000000000000000000 + 
0_10000000110000000000000000000000 = 
1_11000111000000000000000000000000
(4 * w[7])_trunc_3_4 = 111_0001, "belongs to [-Inf, m[-1])" -> q[8] = -2
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
010_1001 + 100_1000 = 111_0001, "belongs to [-Inf, m[-1])" -> q[8] = -2
q_pos = 0000_0000_0001_0000
q_neg = 0000_0000_0000_0110

// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w_sum[8] = csa_sum(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
1_00010010011111111111111111000000
w_carry[8] = csa_carry(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
1_00001011000000000000000001000000
w[8] = w[7] << 2 - q[8] * D = 
1_00011100000000000000000000000000 + 
1_00000001100000000000000000000000 = 
0_00011101100000000000000000000000 >= 0

w_sum[8][(2*WIDTH-1):WIDTH] + w_carry[8][(2*WIDTH-1):WIDTH] = 
0001001001111111 + 
0000101100000000 = 
0001110101111111 = 0001110110000000 - 1

不难发现只要迭代过程中出现过正的商(显然, CLZ_DIFF >= 1时一定会出现)，则最后使用"sum/carry"求出最终余数的时候, 16-bit的Full Adder的"cin = 1".
因此可以使用一个"inc_flag"来记录迭代过程中是否出现过正的商:
for(i = 1; i <= (WIDTH / 2); i++)
	inc_flag = inc_flag | (q[i] >= +1);

于是有:
w[final] = w_sum[final][(2*WIDTH-1):WIDTH] + w_carry[final][(2*WIDTH-1):WIDTH] + inc_flag;

rem = (w[8])_reduced >> CLZ_D = 
0001110110000000 >> 6
0000000001110110

q_final = corr(q_pos - q_neg) = 0000000000001010
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------


// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 24
ITN_W = (2 * WIDTH) + 1 = 49
0_000000000000000000000000000000000000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 100010101001010010010100 = 9082004
D[WIDTH-1:0] = 000100110011001110001001 = 1258377
Q[WIDTH-1:0] = X / D = 7 = 000000000000000000000111
REM[WIDTH-1:0] = 9082004 - 1258377 * 7 = 273365 = 000001000010101111010101

CLZ_X = 0
CLZ_D = 3
CLZ_DIFF = CLZ_D - CLZ_X = 3
Normalized_D = 100110011001110001001000
根据D的值, 可得选择常数:
m[-1] = -14
m[ 0] = - 4
m[+1] = + 4
m[+2] = +14

+ D[ITN_W-1:0] = 0_100110011001110001001000000000000000000000000000
+2D[ITN_W-1:0] = 1_001100110011100010010000000000000000000000000000
- D[ITN_W-1:0] = 1_011001100110001110111000000000000000000000000000
-2D[ITN_W-1:0] = 0_110011001100011101110000000000000000000000000000
~ D[ITN_W-1:0] = 1_011001100110001110110111111111111111111111111111
~2D[ITN_W-1:0] = 0_110011001100011101101111111111111111111111111111

l_shift_num = CLZ_D = 3
shifted_dividend[ITN_W-1:0] = {{0, {(WIDTH){1'b0}}, X[WIDTH-1:0]} << l_shift_num} = 
0_000000000000000000000000100010101001010010010100 << 3 = 
0_000000000000000000000100010101001010010010100000

// ---------------------------------------------------------------------------------------------------------------------------------------
初始化:
w_sum[0][ITN_W-1:0] 	= 0_000000000000000000000100010101001010010010100000
w_carry[0][ITN_W-1:0] 	= 0_000000000000000000000000000000000000000000000000
w[0] 					= 0_000000000000000000000100010101001010010010100000
(4 * w[0])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[1] = 0
q_pos = 00
q_neg = 00

ITER[0]:
w_sum[1] = csa_sum(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_000000000000000000010001010100101001001010000000
w_carry[1] = csa_carry(4 * w_sum[0], 4 * w_carry[0], -q[1] * D) = 
0_000000000000000000000000000000000000000000000000
w[1] = w[0] << 2 - q[1] * D = 
0_000000000000000000010001010100101001001010000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000000000000010001010100101001001010000000
(4 * w[1])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
(4 * w_sum[1])_trunc_3_4 + (4 * w_carry[1])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[2] = 0
q_pos = 0000
q_neg = 0000

ITER[1]:
w_sum[2] = csa_sum(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_000000000000000001000101010010100100101000000000
w_carry[2] = csa_carry(4 * w_sum[1], 4 * w_carry[1], -q[2] * D) = 
0_000000000000000000000000000000000000000000000000
w[2] = w[1] << 2 - q[2] * D = 
0_000000000000000001000101010010100100101000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000000000001000101010010100100101000000000
(4 * w[2])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
(4 * w_sum[2])_trunc_3_4 + (4 * w_carry[2])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[3] = 0
q_pos = 0000_00
q_neg = 0000_00

ITER[2]:
w_sum[3] = csa_sum(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_000000000000000100010101001010010010100000000000
w_carry[3] = csa_carry(4 * w_sum[2], 4 * w_carry[2], -q[3] * D) = 
0_000000000000000000000000000000000000000000000000
w[3] = w[2] << 2 - q[3] * D = 
0_000000000000000100010101001010010010100000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000000000100010101001010010010100000000000
(4 * w[3])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
(4 * w_sum[3])_trunc_3_4 + (4 * w_carry[3])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[4] = 0
q_pos = 0000_0000
q_neg = 0000_0000

ITER[3]:
w_sum[4] = csa_sum(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_000000000000010001010100101001001010000000000000
w_carry[4] = csa_carry(4 * w_sum[3], 4 * w_carry[3], -q[4] * D) = 
0_000000000000000000000000000000000000000000000000
w[4] = w[3] << 2 - q[4] * D = 
0_000000000000010001010100101001001010000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000000010001010100101001001010000000000000
(4 * w[4])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
(4 * w_sum[4])_trunc_3_4 + (4 * w_carry[4])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[5] = 0
q_pos = 0000_0000_00
q_neg = 0000_0000_00

ITER[4]:
w_sum[5] = csa_sum(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
0_000000000001000101010010100100101000000000000000
w_carry[5] = csa_carry(4 * w_sum[4], 4 * w_carry[4], -q[5] * D) = 
0_000000000000000000000000000000000000000000000000
w[5] = w[4] << 2 - q[5] * D = 
0_000000000001000101010010100100101000000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000001000101010010100100101000000000000000
(4 * w[5])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
(4 * w_sum[5])_trunc_3_4 + (4 * w_carry[5])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[6] = 0
q_pos = 0000_0000_0000
q_neg = 0000_0000_0000

ITER[5]:
w_sum[6] = csa_sum(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
0_000000000100010101001010010010100000000000000000
w_carry[6] = csa_carry(4 * w_sum[5], 4 * w_carry[5], -q[6] * D) = 
0_000000000000000000000000000000000000000000000000
w[6] = w[5] << 2 - q[6] * D = 
0_000000000100010101001010010010100000000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000000100010101001010010010100000000000000000
(4 * w[6])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
(4 * w_sum[6])_trunc_3_4 + (4 * w_carry[6])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[7] = 0
q_pos = 0000_0000_0000_00
q_neg = 0000_0000_0000_00

ITER[6]:
w_sum[7] = csa_sum(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
0_000000010001010100101001001010000000000000000000
w_carry[7] = csa_carry(4 * w_sum[6], 4 * w_carry[6], -q[7] * D) = 
0_000000000000000000000000000000000000000000000000
w[7] = w[6] << 2 - q[7] * D = 
0_000000010001010100101001001010000000000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000000010001010100101001001010000000000000000000
(4 * w[7])_trunc_3_4 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
(4 * w_sum[7])_trunc_3_4 + (4 * w_carry[7])_trunc_3_4 = 
000_0000 + 000_0000 = 000_0000, "belongs to [m[0], m[+1])" -> q[8] = 0
q_pos = 0000_0000_0000_0000
q_neg = 0000_0000_0000_0000

ITER[7]:
w_sum[8] = csa_sum(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
0_000001000101010010100100101000000000000000000000
w_carry[8] = csa_carry(4 * w_sum[7], 4 * w_carry[7], -q[8] * D) = 
0_000000000000000000000000000000000000000000000000
w[8] = w[7] << 2 - q[8] * D = 
0_000001000101010010100100101000000000000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000001000101010010100100101000000000000000000000
(4 * w[8])_trunc_3_4 = 000_0001, "belongs to [m[0], m[+1])" -> q[9] = 0
(4 * w_sum[8])_trunc_3_4 + (4 * w_carry[8])_trunc_3_4 = 
000_0001 + 000_0000 = 000_0001, "belongs to [m[0], m[+1])" -> q[9] = 0
q_pos = 0000_0000_0000_0000_00
q_neg = 0000_0000_0000_0000_00

ITER[8]:
w_sum[9] = csa_sum(4 * w_sum[8], 4 * w_carry[8], -q[9] * D) = 
0_000100010101001010010010100000000000000000000000
w_carry[9] = csa_carry(4 * w_sum[8], 4 * w_carry[8], -q[9] * D) = 
0_000000000000000000000000000000000000000000000000
w[9] = w[8] << 2 - q[9] * D = 
0_000100010101001010010010100000000000000000000000 + 
0_000000000000000000000000000000000000000000000000 = 
0_000100010101001010010010100000000000000000000000
(4 * w[9])_trunc_3_4 = 000_0100, "belongs to [m[+1], m[+2])" -> q[10] = +1
(4 * w_sum[9])_trunc_3_4 + (4 * w_carry[9])_trunc_3_4 = 
000_0100 + 000_0000 = 000_0100, "belongs to [m[+1], m[+2])" -> q[10] = +1
q_pos = 0000_0000_0000_0000_0001
q_neg = 0000_0000_0000_0000_0000

ITER[9]:
w_sum[10] = csa_sum(4 * w_sum[9], 4 * w_carry[9], -q[10] * D) = 
1_001000110010100111111101111111111111111111111111
w_carry[10] = csa_carry(4 * w_sum[9], 4 * w_carry[9], -q[10] * D) = 
0_100010001000010000000100000000000000000000000001
w[10] = w[9] << 2 - q[10] * D = 
0_010001010100101001001010000000000000000000000000 + 
1_011001100110001110111000000000000000000000000000 = 
1_101010111010111000000010000000000000000000000000
(4 * w[10])_trunc_3_4 = 110_1010, "belongs to [-Inf, m[-1])" -> q[11] = -2
(4 * w_sum[10])_trunc_3_4 + (4 * w_carry[10])_trunc_3_4 = 
100_1000 + 010_0010 = 110_1010, "belongs to [-Inf, m[-1])" -> q[11] = -2
q_pos = 0000_0000_0000_0000_0001_00
q_neg = 0000_0000_0000_0000_0000_10

ITER[10]:
w_sum[11] = csa_sum(4 * w_sum[10], 4 * w_carry[10], -q[11] * D) = 
1_100111011000111101110111111111111111111111111000
w_carry[11] = csa_carry(4 * w_sum[10], 4 * w_carry[10], -q[11] * D) = 
0_010001000110000100100000000000000000000000001000
w[11] = w[10] << 2 - q[11] * D = 
0_101011101011100000001000000000000000000000000000 + 
1_001100110011100010010000000000000000000000000000 = 
1_111000011111000010011000000000000000000000000000
(4 * w[11])_trunc_3_4 = 111_1000, "belongs to [m[-1], m[0])" -> q[12] = -1
(4 * w_sum[11])_trunc_3_4 + (4 * w_carry[11])_trunc_3_4 = 
110_0111 + 001_0001 = 111_1000, "belongs to [m[-1], m[0])" -> q[12] = -1
q_pos = 0000_0000_0000_0000_0001_0000
q_neg = 0000_0000_0000_0000_0000_1001



// ---------------------------------------------------------------------------------------------------------------------------------------
// 后处理
w_sum[12] = csa_sum(4 * w_sum[11], 4 * w_carry[11], -q[12] * D) = 
1_111111100010010100010111111111111111111111000000
w_carry[12] = csa_carry(4 * w_sum[11], 4 * w_carry[11], -q[12] * D) = 
0_001000110011100110010000000000000000000001000000
w[12] = {w[11] << 2, temp_dividend[11][(WIDTH-1) -: 2]} - q[12] * D = 
1_100001111100001001100000000000000000000000000000 + 
0_100110011001110001001000000000000000000000000000 = 
0_001000010101111010101000000000000000000000000000 >= 0

inc_flag = 1;
w[final] = w_sum[final][(2*WIDTH-1):WIDTH] + w_carry[final][(2*WIDTH-1):WIDTH] + inc_flag = 
111111100010010100010111 + 
001000110011100110010000 + 
1 = 
001000010101111010101000

rem = (w[12])_reduced >> CLZ_D = 
001000010101111010101000 >> 3 = 
000001000010101111010101

q_final = corr(q_pos - q_neg) = 0111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------





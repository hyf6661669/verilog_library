a = 1.00000000000
b = 0.10000010001
a / b = 1.11110111101000111000100011111001110110100010000100
a_scaled = a << 1 = 10.00000000000000
b_scaled = b << 1 = 01.00000100010000

d   = 00100000100010000
2d  = 01000001000100000
~d  = 11011111011101111
~2d = 10111110111011111
-d  = 11011111011110000
-2d = 10111110111100000

// ==================================================================================================
rem_init = 00010000000000000
rem_s[0] = rem_init = 00010000000000000
rem_c[0] = 00000000000000000
rem[0] = 00010000000000000

// ================
// BigIter[0]
d   = 00100000100010000
2d  = 01000001000100000
~d  = 11011111011101111
~2d = 10111110111011111
-d  = 11011111011110000
-2d = 10111110111100000
// ================
// stage[0]
rem_s[0][14:9] + rem_c[0][14:9] = 
010001 + 
000000 = 
010001, belongs to "[13/8, 31/8]" -> q[0] = +2
q_pos = 10
q_neg = 00
q_pos - q_neg = 10
a / b = 1.11110111101000111000100011111001110110100010000100

// stage[1]
rem_s[1] = 01000000000000000
rem_c[1] = 10111110111100000
-> 
rem[1] = 
00010000000000000 + 
11011111011110000 = 
11101111011110000

rem_s[1][14:9] + rem_c[1][14:9] = 
000000 + 
111110 = 
111110, belongs to "[-3/8, 3/8]" -> q[1] = 0
q_pos = 1000
q_neg = 0000
q_pos - q_neg = 1000
a / b = 1.11110111101000111000100011111001110110100010000100

// TODO
adder_9b = (rem_s[1] << 2)[16:8] + (rem_c[1] << 2)[16:8] = 
000000000 + 
111110111 =
000001011
adder_9b[8:3] = 000011, 此时adder_9b[3].carry = 0, 按照TABLE II(b), 应该选择q[1] = +1
->
q_pos = 0101
q_neg = 0000
q_pos - q_neg = 0101
a / b = 1.11110111101000111000100011111001110110100010000100

// stage[2]
rem_s[2] = 11110111010011000
rem_c[2] = 00000001011001000
->
rem[2] = 
10110000110000000 + 
01000111111100000 = 
11111000101100000

rem_s[2][14:9] + rem_c[2][14:9] = 
110111 + 
000001 = 
111000, belongs to "[-12/8, -5/8]" -> q[2] = -1
q_pos = 100000
q_neg = 001001
q_pos - q_neg = 010111
a / b = 1.0111001011111101000110111100110......

adder_7b = ((-q[1] * d) << 2)[16:10] + adder_9b[6:0]
0001111 +
1100001 = 
1110000, adder_7b[6:1] = 111000, belongs to "[-12/8, -4/8]" -> q[2] = -1
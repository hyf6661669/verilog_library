接"test_2.sv", 使用右移的方式:
r_shift_num = log2(N) - 1 - ((CLZ_DIFF) % log2(N));
N =  4 -> r_shift_num = 1 - ((CLZ_DIFF) % 2);
N =  8 -> r_shift_num = 2 - ((CLZ_DIFF) % 3);
N = 16 -> r_shift_num = 3 - ((CLZ_DIFF) % 4);
N = 32 -> r_shift_num = 4 - ((CLZ_DIFF) % 5);
N = 64 -> r_shift_num = 6 - ((CLZ_DIFF) % 6);

// ---------------------------------------------------------------------------------------------------------------------------------------
WIDTH = 28;
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
将3个Radix-2叠加起来形成Radix-8算法, 即:
N = 8;
(WIDTH + 1 + log2(N)) = 32;
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000110100001110011100100011 = 13690659
D[WIDTH-1:0] = 0000000001001001110111011100 = 302556
Q[WIDTH-1:0] = X / D = 45 = 0000000000000000000000101101
REM[WIDTH-1:0] = 13690659 - 302556 * 45 = 75639 = 0000000000010010011101110111

CLZ_X = 4
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 5
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 2 - (5 % 3) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(6 / 3) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1101000011100111001000110000
Divisor[WIDTH-1:0] 		= 1001001110111011100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00100111011101110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_01001110111011100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11011000100010010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_10110001000100100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6] = 000_10010011101110111000000000000 >= 0;
(w[final] / 2) + (-D) = 000_01001001110111011100000000000 + 110_11011000100010010000000000000 = 
11100100010011001101100000000000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1011_01
q_neg = 0000_00

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 101101;
(w[final] / 2) "belongs to [0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 101101;

(w[final] / 2) "belongs to [0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
0010010011101110111000000000 >> 9
0000000000010010011101110111
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_10100001110011100100011000000
w_sum_translation[0] = w_sum[0] =  001_10100001110011100100011000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_01000011100111001000110000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_10110001000100100000000000000
w_sum_translation[1] = 001_01000011100111001000110000000
w_carry_translation[1] = 111_10110001000100100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_11 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_10100001110011100100011000000 +
	110_11011000100010010000000000000
) = 2 * 000_01111010010101110100011000000 = 
000_11110100101011101000110000000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
010_10000111001110010001100000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_01100010001001000000000000000
w_sum_translation[2] = 000_10000111001110010001100000000
w_carry_translation[2] = 001_01100010001001000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_01 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_11110100101011101000110000000 +
	000_00000000000000000000000000000
) = 2 * 000_11110100101011101000110000000 = 
001_11101001010111010001100000000
q_pos = 101
q_neg = 000

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
110_01111011001010000011000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_00001000101001000000000000000
w_sum_translation[3] = 000_01111011001010000011000000000
w_carry_translation[3] = 001_00001000101001000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_01 -> q[4] = +1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_11101001010111010001100000000 +
	110_11011000100010010000000000000
) = 2 * 000_11000001111001100001100000000 = 
001_10000011110011000011000000000
q_pos = 1011
q_neg = 0000

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_01010110000010100110000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_01100010101000000000000000000
w_sum_translation[4] = 111_01010110000010100110000000000
w_carry_translation[4] = 001_01100010101000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_01 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	001_10000011110011000011000000000 +
	110_11011000100010010000000000000
) = 2 * 000_01011100010101010011000000000 = 
000_10111000101010100110000000000
q_pos = 1011_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
110_10101100000101001100000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
010_11000101010000000000000000000
w_sum_translation[5] = 000_10101100000101001100000000000
w_carry_translation[5] = 000_11000101010000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_00 -> q[6] = +1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_10111000101010100110000000000 +
	000_00000000000000000000000000000
) = 2 * 000_10111000101010100110000000000 = 
001_01110001010101001100000000000
q_pos = 1011_01
q_neg = 0000_00

w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	001_01110001010101001100000000000 +
	110_11011000100010010000000000000
) = 2 * 000_01001001110111011100000000000 = 
000_10010011101110111000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000000101000101000011000010 = 1331394
D[WIDTH-1:0] = 0000000000010011100001111111 = 79999
Q[WIDTH-1:0] = X / D = 16 = 0000000000000000000000010000
REM[WIDTH-1:0] = 1331394 - 79999 * 16 = 51410 = 0000000000001100100011010010

CLZ_X = 7
CLZ_D = 11
CLZ_DIFF = CLZ_D - CLZ_X = 4
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 2 - (4 % 3) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(5 / 3) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1010001010000110000100000000
Divisor[WIDTH-1:0] 		= 1001110000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00111000011111110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_01110000111111100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11000111100000010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_10001111000000100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6] = 001_10010001101001000000000000000 >= 0;
(w[final] / 2) + (-D) = 000_11001000110100100000000000000 + 110_11000111100000010000000000000 = 
11110010000010100110000000000000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1000_00
q_neg = 0100_00

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 00010000;
(w[final] / 2) "belongs to [0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 00010000;

(w[final] / 2) "belongs to [0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
0110010001101001000000000000 >> 11
0000000000001100100011010010
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_10100010100001100001000000000
w_sum_translation[0] = w_sum[0] =  000_10100010100001100001000000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
001_01000101000011000010000000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_10001111000000100000000000000
w_sum_translation[1] = 111_01000101000011000010000000000
w_carry_translation[1] = 111_10001111000000100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_10100010100001100001000000000 +
	110_11000111100000010000000000000
) = 2 * 111_01101010000001110001000000000 = 
110_11010100000011100010000000000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_11100100111000100100000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_00110100001110000000000000000
w_sum_translation[2] = 001_11100100111000100100000000000
w_carry_translation[2] = 110_00110100001110000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_11010100000011100010000000000 +
	001_00111000011111110000000000000
) = 2 * 000_00001100100011010010000000000 = 
000_00011001000110100100000000000
q_pos = 100
q_neg = 010

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_11001001110001001000000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_01101000011100000000000000000
w_sum_translation[3] = 001_11001001110001001000000000000
w_carry_translation[3] = 110_01101000011100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_00011001000110100100000000000 +
	000_00000000000000000000000000000
) = 2 * 000_00011001000110100100000000000 = 
000_00110010001101001000000000000
q_pos = 1000
q_neg = 0100

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_10010011100010010000000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_11010000111000000000000000000
w_sum_translation[4] = 001_10010011100010010000000000000
w_carry_translation[4] = 110_11010000111000000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_10 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_00110010001101001000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_00110010001101001000000000000 = 
000_01100100011010010000000000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_00100111000100100000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
101_10100001110000000000000000000
w_sum_translation[5] = 001_00100111000100100000000000000
w_carry_translation[5] = 111_10100001110000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_11 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_01100100011010010000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_01100100011010010000000000000 = 
000_11001000110100100000000000000
q_pos = 1000_00
q_neg = 0100_00

w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_11001000110100100000000000000 +
	000_00000000000000000000000000000
) = 2 * 000_11001000110100100000000000000 = 
001_10010001101001000000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0000001000001011111100000010 = 2146050
D[WIDTH-1:0] = 0000000001000010000111111100 = 270844
Q[WIDTH-1:0] = X / D = 7 = 0000000000000000000000000111
REM[WIDTH-1:0] = 2146050 - 270844 * 7 = 250142 = 0000000000111101000100011110

CLZ_X = 6
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 3
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 2 - (3 % 3) = 2;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(4 / 3) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000001011111100000010000000
Divisor[WIDTH-1:0] 		= 1000010000111111100000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_00001000011111110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_00010000111111100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_11110111100000010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_11101111000000100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[6] = 101_11000110100100110000000000000 < 0;
(w[final] / 2) + (D) = 110_11100011010010011000000000000 + 001_00001000011111110000000000000 = 
11111101011110010001000000000000 < 0 -> (w[final] / 2) "belongs to [-2D, -D)";
// 最后一次迭代的商
q_pos = 1000_00
q_neg = 0101_11

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 1001;
(w[final] / 2) "belongs to [-2D, -D)" -> quotient_correction_coefficient = -2;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 0111;

(w[final] / 2) "belongs to [-2D, -D)" -> remainder_correction_coefficient = -2;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
(110_11100011010010011000000000000 + 010_00010000111111100000000000000) >> 9 = 
0111101000100011110000000000 >> 9
0000000000111101000100011110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_01000001011111100000010000000
w_sum_translation[0] = w_sum[0] =  000_01000001011111100000010000000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_00000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_10000010111111000000100000000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_11101111000000100000000000000
w_sum_translation[1] = 110_10000010111111000000100000000
w_carry_translation[1] = 111_11101111000000100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_01000001011111100000010000000 +
	110_11110111100000010000000000000
) = 2 * 111_00111000111111110000010000000 = 
110_01110001111111100000100000000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_11001011000000100001000000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_00101001111110000000000000000
w_sum_translation[2] = 000_11001011000000100001000000000
w_carry_translation[2] = 110_00101001111110000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_01110001111111100000100000000 +
	001_00001000011111110000000000000
) = 2 * 111_01111010011111010000100000000 = 
110_11110100111110100001000000000
q_pos = 100
q_neg = 010

// 第2次大迭代
w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
001_10010110000001000010000000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_01010011111100000000000000000
w_sum_translation[3] = 111_10010110000001000010000000000
w_carry_translation[3] = 110_01010011111100000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_10 -> q[4] = -1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	110_11110100111110100001000000000 +
	000_00000000000000000000000000000
) = 2 * 110_11110100111110100001000000000 = 
101_11101001111101000010000000000
q_pos = 1000
q_neg = 0101

w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_10011011000101100100000000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_01001001110100000000000000000
w_sum_translation[4] = 111_10011011000101100100000000000
w_carry_translation[4] = 110_01001001110100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_10 -> q[5] = -1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	101_11101001111101000010000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11110010011100110010000000000 = 
101_11100100111001100100000000000
q_pos = 1000_0
q_neg = 0101_1

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
001_10110101011100101000000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
100_00100101010110000000000000000
w_sum_translation[5] = 111_10110101011100101000000000000
w_carry_translation[5] = 110_00100101010110000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 11_10 -> q[6] = -1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	101_11100100111001100100000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11101101011001010100000000000 = 
101_11011010110010101000000000000
q_pos = 1000_00
q_neg = 0101_11


w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	101_11011010110010101000000000000 +
	001_00001000011111110000000000000
) = 2 * 110_11100011010010011000000000000 = 
101_11000110100100110000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
// ---------------------------------------------------------------------------------------------------------------------------------------
将4个Radix-2叠加起来形成Radix-16算法, 即:
N = 16;
(WIDTH + 1 + log2(N)) = 33;
// ---------------------------------------------------------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 0111111111100010111011110011 = 134098675
D[WIDTH-1:0] = 0000000011110001000101000011 = 987459
Q[WIDTH-1:0] = X / D = 135 = 0000000000000000000010000111
REM[WIDTH-1:0] = 134098675 - 987459 * 135 = 791710 = 0000000011000001010010011110

CLZ_X = 1
CLZ_D = 8
CLZ_DIFF = CLZ_D - CLZ_X = 7
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (7 % 4) = 0;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(8 / 4) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111111111000101110111100110
Divisor[WIDTH-1:0] 		= 1111000100010100001100000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_111000100010100001100000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 011_110001000101000011000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_000111011101011110100000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 100_001110111010111101000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8] = 011_000001010010011110000000000000 >= 0;
(w[final] / 2) + (-D) = 001_100000101001001111000000000000 + 110_000111011101011110100000000000 = 
111_101000000110101101100000000000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1000_1000
q_neg = 0000_0001

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 10000111;
(w[final] / 2) "belongs to [0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 10000111;

(w[final] / 2) "belongs to [0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
1100000101001001111000000000 >> 8 =
0000000011000001010010011110
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  001_111111111000101110111100110000
w_sum_translation[0] = w_sum[0] =  001_111111111000101110111100110000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 01_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
011_111111110001011101111001100000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_001110111010111101000000000000
w_sum_translation[1] = 001_111111110001011101111001100000
w_carry_translation[1] = 110_001110111010111101000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 01_10 -> q[2] = 0
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	001_111111111000101110111100110000 +
	110_000111011101011110100000000000
) = 2 * 000_000111010110001101011100110000 = 
000_001110101100011010111001100000
q_pos = 10
q_neg = 00

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
011_111111100010111011110011000000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
100_011101110101111010000000000000
w_sum_translation[2] = 001_111111100010111011110011000000
w_carry_translation[2] = 110_011101110101111010000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 01_10 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	000_001110101100011010111001100000 +
	000_000000000000000000000000000000
) = 2 * 000_001110101100011010111001100000 = 
000_011101011000110101110011000000
q_pos = 100
q_neg = 000

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
011_111111000101110111100110000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_111011101011110100000000000000
w_sum_translation[3] = 001_111111000101110111100110000000
w_carry_translation[3] = 110_111011101011110100000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 01_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_011101011000110101110011000000 +
	000_000000000000000000000000000000
) = 2 * 000_011101011000110101110011000000 = 
000_111010110001101011100110000000
q_pos = 1000
q_neg = 0000

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
011_111110001011101111001100000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
101_110111010111101000000000000000
w_sum_translation[4] = 001_111110001011101111001100000000
w_carry_translation[4] = 111_110111010111101000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 01_11 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_111010110001101011100110000000 +
	000_000000000000000000000000000000
) = 2 * 000_111010110001101011100110000000 = 
001_110101100011010111001100000000
q_pos = 1000_0
q_neg = 0000_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
011_111100010111011110011000000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_101110101111010000000000000000
w_sum_translation[5] = 001_111100010111011110011000000000
w_carry_translation[5] = 001_101110101111010000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 01_01 -> q[6] = +2
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	001_110101100011010111001100000000 +
	000_000000000000000000000000000000
) = 2 * 001_110101100011010111001100000000 = 
011_101011000110101110011000000000
q_pos = 1000_10
q_neg = 0000_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
100_111000000101100110110000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_111011111101110000000000000000
w_sum_translation[6] = 110_111000000101100110110000000000
w_carry_translation[6] = 000_111011111101110000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 10_00 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	011_101011000110101110011000000000 +
	100_001110111010111101000000000000
) = 2 * 111_111010000001101011011000000000 = 
111_110100000011010110110000000000
q_pos = 1000_100
q_neg = 0000_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
101_110000001011001101100000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
001_110111111011100000000000000000
w_sum_translation[7] = 111_110000001011001101100000000000
w_carry_translation[7] = 111_110111111011100000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 11_11 -> q[8] = -1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	111_110100000011010110110000000000 +
	000_000000000000000000000000000000
) = 2 * 111_110100000011010110110000000000 = 
111_101000000110101101100000000000
q_pos = 1000_1000
q_neg = 0000_0001

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	111_101000000110101101100000000000 +
	001_111000100010100001100000000000
) = 2 * 001_100000101001001111000000000000 = 
011_000001010010011110000000000000



// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1111111111100010111011110011 = 268316403
D[WIDTH-1:0] = 0000000000111111000101001111 = 258383
Q[WIDTH-1:0] = X / D = 1038 = 0000000000000000010000001110
REM[WIDTH-1:0] = 268316403 - 258383 * 1038 = 114849 = 0000000000011100000010100001

CLZ_X = 0
CLZ_D = 10
CLZ_DIFF = CLZ_D - CLZ_X = 10
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (10 % 4) = 1;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(11 / 4) = 3;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1111111111100010111011110011
Divisor[WIDTH-1:0] 		= 1111110001010011110000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_111110001010011110000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 011_111100010100111100000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_000001110101100010000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 100_000011101011000100000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[12] = 001_110000001010000100000000000000 >= 0;
(w[final] / 2) + (-D) = 000_111000000101000010000000000000 + 110_000111011101011110100000000000 = 
110_111111100010100000100000000000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1000_0001_0000
q_neg = 0100_0000_0010

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 010000001110;
(w[final] / 2) "belongs to [0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 010000001110;

(w[final] / 2) "belongs to [0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
0111000000101000010000000000 >> 10 =
0000000000011100000010100001
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_111111111110001011101111001100
w_sum_translation[0] = w_sum[0] =  000_111111111110001011101111001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
001_111111111100010111011110011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_000011101011000100000000000000
w_sum_translation[1] = 111_111111111100010111011110011000
w_carry_translation[1] = 110_000011101011000100000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 11_10 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_111111111110001011101111001100 +
	110_000001110101100010000000000000
) = 2 * 111_000001110011101101101111001100 = 
110_000011100111011011011110011000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
000_000100111010011010111100110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
111_111110101001011000000000000000
w_sum_translation[2] = 000_000100111010011010111100110000
w_carry_translation[2] = 111_111110101001011000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_11 -> q[3] = 0
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_000011100111011011011110011000 +
	001_111110001010011110000000000000
) = 2 * 000_000001110001111001011110011000 = 
000_000011100011110010111100110000
q_pos = 100
q_neg = 010

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
000_001001110100110101111001100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
111_111101010010110000000000000000
w_sum_translation[3] = 000_001001110100110101111001100000
w_carry_translation[3] = 111_111101010010110000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_11 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	000_000011100011110010111100110000 +
	000_000000000000000000000000000000
) = 2 * 000_000011100011110010111100110000 = 
000_000111000111100101111001100000
q_pos = 1000
q_neg = 0100

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
000_010011101001101011110011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
111_111010100101100000000000000000
w_sum_translation[4] = 000_010011101001101011110011000000
w_carry_translation[4] = 111_111010100101100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_11 -> q[5] = 0
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	000_000111000111100101111001100000 +
	000_000000000000000000000000000000
) = 2 * 000_000111000111100101111001100000 = 
000_001110001111001011110011000000
q_pos = 1000_0
q_neg = 0100_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_100111010011010111100110000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
111_110101001011000000000000000000
w_sum_translation[5] = 000_100111010011010111100110000000
w_carry_translation[5] = 111_110101001011000000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 00_11 -> q[6] = 0
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	000_001110001111001011110011000000 +
	000_000000000000000000000000000000
) = 2 * 000_001110001111001011110011000000 = 
000_011100011110010111100110000000
q_pos = 1000_00
q_neg = 0100_00

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
001_001110100110101111001100000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
111_101010010110000000000000000000
w_sum_translation[6] = 001_001110100110101111001100000000
w_carry_translation[6] = 111_101010010110000000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 01_11 -> q[7] = 0
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	000_011100011110010111100110000000 +
	000_000000000000000000000000000000
) = 2 * 000_011100011110010111100110000000 = 
000_111000111100101111001100000000
q_pos = 1000_000
q_neg = 0100_000

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
010_011101001101011110011000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
111_010100101100000000000000000000
w_sum_translation[7] = 000_011101001101011110011000000000
w_carry_translation[7] = 001_010100101100000000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 00_01 -> q[8] = +1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	000_111000111100101111001100000000 +
	000_000000000000000000000000000000
) = 2 * 000_111000111100101111001100000000 = 
001_110001111001011110011000000000
q_pos = 1000_0001
q_neg = 0100_0000

// 第3次大迭代
w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
110_010000101001111000110000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
001_010110110100001000000000000000
w_sum_translation[8] = 110_010000101001111000110000000000
w_carry_translation[8] = 001_010110110100001000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 10_01 -> q[9] = 0
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	001_110001111001011110011000000000 +
	110_000001110101100010000000000000
) = 2 * 111_110011101111000000011000000000 = 
111_100111011110000000110000000000
q_pos = 1000_0001_0
q_neg = 0100_0000_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
100_100001010011110001100000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
010_101101101000010000000000000000
w_sum_translation[9] = 110_100001010011110001100000000000
w_carry_translation[9] = 000_101101101000010000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_00 -> q[10] = 0
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	111_100111011110000000110000000000 +
	000_000000000000000000000000000000
) = 2 * 111_100111011110000000110000000000 = 
111_001110111100000001100000000000
q_pos = 1000_0001_00
q_neg = 0100_0000_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
101_000010100111100011000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_011011010000100000000000000000
w_sum_translation[10] = 111_000010100111100011000000000000
w_carry_translation[10] = 111_011011010000100000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 11_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	111_001110111100000001100000000000 +
	000_000000000000000000000000000000
) = 2 * 111_001110111100000001100000000000 = 
110_011101111000000011000000000000
q_pos = 1000_0001_000
q_neg = 0100_0000_001

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
011_001111111010111010000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
101_101000001010001000000000000000
w_sum_translation[11] = 001_001111111010111010000000000000
w_carry_translation[11] = 111_101000001010001000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 01_11 -> q[12] = 0
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	110_011101111000000011000000000000 +
	001_111110001010011110000000000000
) = 2 * 000_011100000010100001000000000000 = 
000_111000000101000010000000000000
q_pos = 1000_0001_0000
q_neg = 0100_0000_0010

w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	000_111000000101000010000000000000 +
	000_000000000000000000000000000000
) = 2 * 000_111000000101000010000000000000 = 
001_110000001010000100000000000000




// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1000001000100010111111111100 = 136458236
D[WIDTH-1:0] = 0000000001100001000101001000 = 397640
Q[WIDTH-1:0] = X / D = 343 = 0000000000000000000101010111
REM[WIDTH-1:0] = 136458236 - 397640 * 343 = 67716 = 0000000000010000100010000100

CLZ_X = 0
CLZ_D = 9
CLZ_DIFF = CLZ_D - CLZ_X = 9
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (9 % 4) = 2;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(10 / 4) = 3;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000001000100010111111111100
Divisor[WIDTH-1:0] 		= 1100001000101001000000000000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_100001000101001000000000000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 011_000010001010010000000000000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_011110111010111000000000000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 100_111101110101110000000000000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[12] = 000_100001000100001000000000000000 >= 0;
(w[final] / 2) + (-D) = 000_010000100010000100000000000000 + 110_011110111010111000000000000000 = 
110101111011100111100000000000000 < 0 -> (w[final] / 2) "belongs to [0, +D)";
// 最后一次迭代的商
q_pos = 1010_1010_1001
q_neg = 1001_0101_0010

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 000101010111;
(w[final] / 2) "belongs to [0, +D)" -> quotient_correction_coefficient = 0;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 000101010111;

(w[final] / 2) "belongs to [0, +D)" -> remainder_correction_coefficient = 0;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
0010000100010000100000000000 >> 9 =
0000000000010000100010000100
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_010000010001000101111111111000
w_sum_translation[0] = w_sum[0] =  000_010000010001000101111111111000
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_100000100010001011111111110000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
100_111101110101110000000000000000
w_sum_translation[1] = 110_100000100010001011111111110000
w_carry_translation[1] = 110_111101110101110000000000000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_10 -> q[2] = -2
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_010000010001000101111111111000 +
	110_011110111010111000000000000000
) = 2 * 110_101111001011111101111111111000 = 
101_011110010111111011111111110000
q_pos = 10
q_neg = 10

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
010_111110111011010111111111100000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
110_000010001001000000000000000000
w_sum_translation[2] = 000_111110111011010111111111100000
w_carry_translation[2] = 000_000010001001000000000000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 00_00 -> q[3] = +1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	101_011110010111111011111111110000 +
	011_000010001010010000000000000000
) = 2 * 000_100000100010001011111111110000 = 
001_000001000100010111111111100000
q_pos = 101
q_neg = 100

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
101_000100010001011111111111000000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
001_111011101101000000000000000000
w_sum_translation[3] = 111_000100010001011111111111000000
w_carry_translation[3] = 111_111011101101000000000000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 11_11 -> q[4] = -1
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	001_000001000100010111111111100000 +
	110_011110111010111000000000000000
) = 2 * 111_011111111111001111111111100000 = 
110_111111111110011111111111000000
q_pos = 1010
q_neg = 1001

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
010_111101110010101111111110000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
110_000100010100100000000000000000
w_sum_translation[4] = 000_111101110010101111111110000000
w_carry_translation[4] = 000_000100010100100000000000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 00_00 -> q[5] = +1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	110_111111111110011111111111000000 +
	001_100001000101001000000000000000
) = 2 * 000_100001000011100111111111000000 = 
001_000010000111001111111110000000
q_pos = 1010_1
q_neg = 1001_0

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
101_001110111001101111111100000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
001_110011001010100000000000000000
w_sum_translation[5] = 111_001110111001101111111100000000
w_carry_translation[5] = 111_110011001010100000000000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 11_11 -> q[6] = -1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	001_000010000111001111111110000000 +
	110_011110111010111000000000000000
) = 2 * 111_100001000010000111111110000000 = 
111_000010000100001111111100000000
q_pos = 1010_10
q_neg = 1001_01

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
010_111001101100001111111000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
110_001100100110100000000000000000
w_sum_translation[6] = 000_111001101100001111111000000000
w_carry_translation[6] = 000_001100100110100000000000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 00_00 -> q[7] = +1
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	111_000010000100001111111100000000 +
	001_100001000101001000000000000000
) = 2 * 000_100011001001010111111100000000 = 
001_000110010010101111111000000000
q_pos = 1010_101
q_neg = 1001_010

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
101_010111100000101111110000000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
001_110010111010100000000000000000
w_sum_translation[7] = 111_010111100000101111110000000000
w_carry_translation[7] = 111_110010111010100000000000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 11_11 -> q[8] = -1
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	001_000110010010101111111000000000 +
	110_011110111010111000000000000000
) = 2 * 111_100101001101100111111000000000 = 
111_001010011011001111110000000000
q_pos = 1010_1010
q_neg = 1001_0101

// 第3次大迭代
w_sum[8] = 2 * csa_sum(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
010_001000111110001111100000000000
w_carry[8] = 2 * csa_carry(w_sum_translation[7], w_carry_translation[7], -q[8] * D) = 
111_001110000010100000000000000000
w_sum_translation[8] = 000_001000111110001111100000000000
w_carry_translation[8] = 001_001110000010100000000000000000
{w_sum_translation[8][MSB-1:MSB-2], w_carry_translation[8][MSB-1:MSB-2]} = 00_01 -> q[9] = +1
w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	111_001010011011001111110000000000 +
	001_100001000101001000000000000000
) = 2 * 000_101011100000010111110000000000 = 
001_010111000000101111100000000000
q_pos = 1010_1010_1
q_neg = 1001_0101_0

w_sum[9] = 2 * csa_sum(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
110_110000001100101111000000000000
w_carry[9] = 2 * csa_carry(w_sum_translation[8], w_carry_translation[8], -q[9] * D) = 
000_111011101010100000000000000000
w_sum_translation[9] = 110_110000001100101111000000000000
w_carry_translation[9] = 000_111011101010100000000000000000
{w_sum_translation[9][MSB-1:MSB-2], w_carry_translation[9][MSB-1:MSB-2]} = 10_00 -> q[10] = 0
w[9] = 2 * (w[8] - q[9] * D) = 2 * (
	001_010111000000101111100000000000 +
	110_011110111010111000000000000000
) = 2 * 111_110101111011100111100000000000 = 
111_101011110111001111000000000000
q_pos = 1010_1010_10
q_neg = 1001_0101_00

w_sum[10] = 2 * csa_sum(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
101_100000011001011110000000000000
w_carry[10] = 2 * csa_carry(w_sum_translation[9], w_carry_translation[9], -q[10] * D) = 
001_110111010101000000000000000000
w_sum_translation[10] = 111_100000011001011110000000000000
w_carry_translation[10] = 111_110111010101000000000000000000
{w_sum_translation[10][MSB-1:MSB-2], w_carry_translation[10][MSB-1:MSB-2]} = 11_11 -> q[11] = -1
w[10] = 2 * (w[9] - q[10] * D) = 2 * (
	111_101011110111001111000000000000 +
	000_000000000000000000000000000000
) = 2 * 111_101011110111001111000000000000 = 
111_010111101110011110000000000000
q_pos = 1010_1010_100
q_neg = 1001_0101_001

w_sum[11] = 2 * csa_sum(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
011_101100010010101100000000000000
w_carry[11] = 2 * csa_carry(w_sum_translation[10], w_carry_translation[10], -q[11] * D) = 
110_000101010100100000000000000000
w_sum_translation[11] = 001_101100010010101100000000000000
w_carry_translation[11] = 000_000101010100100000000000000000
{w_sum_translation[11][MSB-1:MSB-2], w_carry_translation[11][MSB-1:MSB-2]} = 01_00 -> q[12] = +1
w[11] = 2 * (w[10] - q[11] * D) = 2 * (
	111_010111101110011110000000000000 +
	001_100001000101001000000000000000
) = 2 * 000_111000110011100110000000000000 = 
001_110001100111001100000000000000
q_pos = 1010_1010_1001
q_neg = 1001_0101_0010

w[12] = 2 * (w[11] - q[12] * D) = 2 * (
	001_110001100111001100000000000000 +
	110_011110111010111000000000000000
) = 2 * 000_010000100010000100000000000000 = 
000_100001000100001000000000000000


// ---------------------------------------------------------------------------------------------------------------------------------------
X[WIDTH-1:0] = 1000010000100010111000001100 = 138554892
D[WIDTH-1:0] = 0000100001111110110101111111 = 8908159
Q[WIDTH-1:0] = X / D = 15 = 0000000000000000000000001111
REM[WIDTH-1:0] = 138554892 - 8908159 * 15 = 4932507 = 0000010010110100001110011011

CLZ_X = 0
CLZ_D = 4
CLZ_DIFF = CLZ_D - CLZ_X = 4
r_shift_num = log2(N) - 1 - (CLZ_DIFF % log2(N)) = 3 - (4 % 4) = 3;
迭代次数
iter_num = ceil((CLZ_DIFF + 1) / log2(N)) = ceil(5 / 4) = 2;
规格化操作之后:
Dividend[WIDTH-1:0] 	= 1000010000100010111000001100
Divisor[WIDTH-1:0] 		= 1000011111101101011111110000

+ D[(WIDTH + 1 + log2(N))-1:0] = 001_000011111101101011111110000000
+2D[(WIDTH + 1 + log2(N))-1:0] = 010_000111111011010111111100000000
- D[(WIDTH + 1 + log2(N))-1:0] = 110_111100000010010100000010000000
-2D[(WIDTH + 1 + log2(N))-1:0] = 101_111000000100101000000100000000
// ---------------------------------------------------------------------------------------------------------------------------------------
// 根据迭代结果计算商和余数
// 最后一次迭代的余数
w[final] = w[8] = 111_000011010101100001110000000000 < 0;
(w[final] / 2) + (D) = 111_100001101010110000111000000000 + 001_000011111101101011111110000000 = 
000_100101101000011100110110000000 >= 0 -> (w[final] / 2) "belongs to [-D, 0)";
// 最后一次迭代的商
q_pos = 1000_0000
q_neg = 0111_0000

q_calculated_pre[WIDTH-1:0] = q_pos[WIDTH-1:0] - q_neg[WIDTH-1:0] = 00010000;
(w[final] / 2) "belongs to [-D, 0)" -> quotient_correction_coefficient = 1;
q_calculated[WIDTH-1:0] = q_calculated_pre[WIDTH-1:0] + quotient_correction_coefficient = 1111;

(w[final] / 2) "belongs to [-D, 0)" -> remainder_correction_coefficient = 1;
remainder_calculated[WIDTH-1:0] = (((w[final] / 2) - remainder_correction_coefficient * D)[(log2(N) - 1) +: WIDTH]) >> CLZ_D = 
(111_100001101010110000111000000000 + 001_000011111101101011111110000000) >> 4 =
0100101101000011100110110000 >> 4 = 
0000010010110100001110011011
// 结果正确
// ---------------------------------------------------------------------------------------------------------------------------------------

初始化:
w[0][(WIDTH + 1 + log2(N))-1:0] =  000_001000010000100010111000001100
w_sum_translation[0] = w_sum[0] =  000_001000010000100010111000001100
w_carry_translation[0] = w_carry[0] = {(WIDTH + 1 + log2(N)){1'b0}} = 000_000000000000000000000000000000
// 第1次大迭代
{w_sum_translation[0][MSB-1:MSB-2], w_carry_translation[0][MSB-1:MSB-2]} = 00_00 -> q[1] = +1
q_pos = 1
q_neg = 0

w_sum[1] = 2 * csa_sum(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
000_010000100001000101110000011000
w_carry[1] = 2 * csa_carry(w_sum_translation[0], w_carry_translation[0], -q[1] * D) = 
101_111000000100101000000100000000
w_sum_translation[1] = 110_010000100001000101110000011000
w_carry_translation[1] = 111_111000000100101000000100000000
{w_sum_translation[1][MSB-1:MSB-2], w_carry_translation[1][MSB-1:MSB-2]} = 10_11 -> q[2] = -1
w[1] = 2 * (w[0] - q[1] * D) = 2 * (
	000_001000010000100010111000001100 +
	110_111100000010010100000010000000
) = 2 * 111_000100010010110110111010001100 = 
110_001000100101101101110100011000
q_pos = 10
q_neg = 01

w_sum[2] = 2 * csa_sum(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
001_010110110000001100010100110000
w_carry[2] = 2 * csa_carry(w_sum_translation[1], w_carry_translation[1], -q[2] * D) = 
101_000010010110100111010000000000
w_sum_translation[2] = 111_010110110000001100010100110000
w_carry_translation[2] = 111_000010010110100111010000000000
{w_sum_translation[2][MSB-1:MSB-2], w_carry_translation[2][MSB-1:MSB-2]} = 11_11 -> q[3] = -1
w[2] = 2 * (w[1] - q[2] * D) = 2 * (
	110_001000100101101101110100011000 +
	001_000011111101101011111110000000
) = 2 * 111_001100100011011001110010011000 = 
110_011001000110110011100100110000
q_pos = 100
q_neg = 011

w_sum[3] = 2 * csa_sum(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
010_101110110110000001110101100000
w_carry[3] = 2 * csa_carry(w_sum_translation[2], w_carry_translation[2], -q[3] * D) = 
100_001011010010111101010000000000
w_sum_translation[3] = 000_101110110110000001110101100000
w_carry_translation[3] = 110_001011010010111101010000000000
{w_sum_translation[3][MSB-1:MSB-2], w_carry_translation[3][MSB-1:MSB-2]} = 00_10 -> q[4] = 0
w[3] = 2 * (w[2] - q[3] * D) = 2 * (
	110_011001000110110011100100110000 +
	001_000011111101101011111110000000
) = 2 * 111_011101000100011111100010110000 = 
110_111010001000111111000101100000
q_pos = 1000
q_neg = 0110

// 第2次大迭代
w_sum[4] = 2 * csa_sum(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
001_011101101100000011101011000000
w_carry[4] = 2 * csa_carry(w_sum_translation[3], w_carry_translation[3], -q[4] * D) = 
100_010110100101111010100000000000
w_sum_translation[4] = 111_011101101100000011101011000000
w_carry_translation[4] = 110_010110100101111010100000000000
{w_sum_translation[4][MSB-1:MSB-2], w_carry_translation[4][MSB-1:MSB-2]} = 11_10 -> q[5] = -1
w[4] = 2 * (w[3] - q[4] * D) = 2 * (
	110_111010001000111111000101100000 +
	000_000000000000000000000000000000
) = 2 * 110_111010001000111111000101100000 = 
101_110100010001111110001011000000
q_pos = 1000_0
q_neg = 0110_1

w_sum[5] = 2 * csa_sum(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
000_010001101000100101101010000000
w_carry[5] = 2 * csa_carry(w_sum_translation[4], w_carry_translation[4], -q[5] * D) = 
101_011110110110101110101000000000
w_sum_translation[5] = 110_010001101000100101101010000000
w_carry_translation[5] = 111_011110110110101110101000000000
{w_sum_translation[5][MSB-1:MSB-2], w_carry_translation[5][MSB-1:MSB-2]} = 10_11 -> q[6] = -1
w[5] = 2 * (w[4] - q[5] * D) = 2 * (
	101_110100010001111110001011000000 +
	001_000011111101101011111110000000
) = 2 * 110_111000001111101010001001000000 = 
101_110000011111010100010010000000
q_pos = 1000_00
q_neg = 0110_11

w_sum[6] = 2 * csa_sum(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
000_011001000111000001111000000000
w_carry[6] = 2 * csa_carry(w_sum_translation[5], w_carry_translation[5], -q[6] * D) = 
101_001111110010111110101000000000
w_sum_translation[6] = 110_011001000111000001111000000000
w_carry_translation[6] = 111_001111110010111110101000000000
{w_sum_translation[6][MSB-1:MSB-2], w_carry_translation[6][MSB-1:MSB-2]} = 10_11 -> q[7] = -1
w[6] = 2 * (w[5] - q[6] * D) = 2 * (
	101_110000011111010100010010000000 +
	001_000011111101101011111110000000
) = 2 * 110_110100011101000000010000000000 = 
101_101000111010000000100000000000
q_pos = 1000_000
q_neg = 0110_111

w_sum[7] = 2 * csa_sum(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
000_101010010000101001011100000000
w_carry[7] = 2 * csa_carry(w_sum_translation[6], w_carry_translation[6], -q[7] * D) = 
100_101111011110101111100000000000
w_sum_translation[7] = 110_101010010000101001011100000000
w_carry_translation[7] = 110_101111011110101111100000000000
{w_sum_translation[7][MSB-1:MSB-2], w_carry_translation[7][MSB-1:MSB-2]} = 10_10 -> q[8] = -2
w[7] = 2 * (w[6] - q[7] * D) = 2 * (
	101_101000111010000000100000000000 +
	001_000011111101101011111110000000
) = 2 * 110_101100110111101100011110000000 = 
101_011001101111011000111100000000
q_pos = 1000_0000
q_neg = 0111_0000

w[8] = 2 * (w[7] - q[8] * D) = 2 * (
	101_011001101111011000111100000000 +
	010_000111111011010111111100000000
) = 2 * 111_100001101010110000111000000000 = 
111_000011010101100001110000000000


